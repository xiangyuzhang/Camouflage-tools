
module c432 (N1, N2, N3, N4, NO);

input N1,N2,N3,N4;

output NO;

wire ;

nand4 gate1( .a(N1), .a(N2), .a(N3), .a(N4), .O(NO) );


endmodule