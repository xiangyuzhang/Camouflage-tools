
module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);

input  N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,CONST1,CONST0 //RE__PI;

input D_0,D_1,D_2,D_3,D_4,D_5,D_6,D_7,D_8,D_9,D_10,D_11,D_12,D_13,D_14,D_15,D_16,D_17,D_18,D_19,D_20,D_21,D_22,D_23,D_24,D_25,D_26,D_27,D_28,D_29,D_30,D_31,D_32,D_33,D_34,D_35,D_36,D_37,D_38,D_39,D_40,D_41 //RE__ALLOW(00,01,10,11);

output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877,D_0_NOT,D_1_NOT,N255_NOT,N255_OBF,ED_0,ED_1,ED_2,ED_3,ED_4,ED_5,ED_6,ED_7,ED_8,ED_9,D_2_NOT,D_3_NOT,N600_NOT,N600_OBF,ED_10,ED_11,ED_12,ED_13,ED_14,ED_15,ED_16,ED_17,ED_18,ED_19,D_4_NOT,D_5_NOT,N739_NOT,N739_OBF,ED_20,ED_21,ED_22,ED_23,ED_24,ED_25,ED_26,ED_27,ED_28,ED_29,D_6_NOT,D_7_NOT,N376_NOT,N376_OBF,ED_30,ED_31,ED_32,ED_33,ED_34,ED_35,ED_36,ED_37,ED_38,ED_39,D_8_NOT,D_9_NOT,N533_NOT,N533_OBF,ED_40,ED_41,ED_42,ED_43,ED_44,ED_45,ED_46,ED_47,ED_48,ED_49,D_10_NOT,D_11_NOT,N451_NOT,N451_OBF,ED_50,ED_51,ED_52,ED_53,ED_54,ED_55,ED_56,ED_57,ED_58,ED_59,D_12_NOT,D_13_NOT,N644_NOT,N644_OBF,ED_60,ED_61,ED_62,ED_63,ED_64,ED_65,ED_66,ED_67,ED_68,ED_69,D_14_NOT,D_15_NOT,N759_NOT,N759_OBF,ED_70,ED_71,ED_72,ED_73,ED_74,ED_75,ED_76,ED_77,ED_78,ED_79,D_16_NOT,D_17_NOT,N17_NOT,N17_OBF,ED_80,ED_81,ED_82,ED_83,ED_84,ED_85,ED_86,ED_87,ED_88,ED_89,D_18_NOT,D_19_NOT,N29_NOT,N29_OBF,ED_90,ED_91,ED_92,ED_93,ED_94,ED_95,ED_96,ED_97,ED_98,ED_99,D_20_NOT,D_21_NOT,N219_NOT,N219_OBF,ED_100,ED_101,ED_102,ED_103,ED_104,ED_105,ED_106,ED_107,ED_108,ED_109,D_22_NOT,D_23_NOT,N130_NOT,N130_OBF,ED_110,ED_111,ED_112,ED_113,ED_114,ED_115,ED_116,ED_117,ED_118,ED_119,D_24_NOT,D_25_NOT,N736_NOT,N736_OBF,ED_120,ED_121,ED_122,ED_123,ED_124,ED_125,ED_126,ED_127,ED_128,ED_129,D_26_NOT,D_27_NOT,N451_NOT,N451_OBF,ED_130,ED_131,ED_132,ED_133,ED_134,ED_135,ED_136,ED_137,ED_138,ED_139,D_28_NOT,D_29_NOT,N228_NOT,N228_OBF,ED_140,ED_141,ED_142,ED_143,ED_144,ED_145,ED_146,ED_147,ED_148,ED_149,D_30_NOT,D_31_NOT,N349_NOT,N349_OBF,ED_150,ED_151,ED_152,ED_153,ED_154,ED_155,ED_156,ED_157,ED_158,ED_159,D_32_NOT,D_33_NOT,N417_NOT,N417_OBF,ED_160,ED_161,ED_162,ED_163,ED_164,ED_165,ED_166,ED_167,ED_168,ED_169,D_34_NOT,D_35_NOT,N830_NOT,N830_OBF,ED_170,ED_171,ED_172,ED_173,ED_174,ED_175,ED_176,ED_177,ED_178,ED_179,D_36_NOT,D_37_NOT,N29_NOT,N29_OBF,ED_180,ED_181,ED_182,ED_183,ED_184,ED_185,ED_186,ED_187,ED_188,ED_189,D_38_NOT,D_39_NOT,N59_NOT,N59_OBF,ED_190,ED_191,ED_192,ED_193,ED_194,ED_195,ED_196,ED_197,ED_198,ED_199,D_40_NOT,D_41_NOT,N557_NOT,N557_OBF,ED_200,ED_201,ED_202,ED_203,ED_204,ED_205,ED_206,ED_207,ED_208,ED_209;


nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );
nand2 gate8( .a(N29), .b(N68), .O(N285) );
nand3 gate9( .a(N59_OBF), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29_OBF), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29_OBF), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );
nand2 gate20( .a(N91), .b(N96), .O(N301) );
or2 gate21( .a(N91), .b(N96), .O(N302) );
nand2 gate22( .a(N101), .b(N106), .O(N303) );
or2 gate23( .a(N101), .b(N106), .O(N304) );
nand2 gate24( .a(N111), .b(N116), .O(N305) );
or2 gate25( .a(N111), .b(N116), .O(N306) );
nand2 gate26( .a(N121), .b(N126), .O(N307) );
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
and2 gate31( .a(N17), .b(N138), .O(N317) );
and2 gate32( .a(N152), .b(N138), .O(N318) );
nand2 gate33( .a(N59), .b(N156), .O(N319) );
nor2 gate34( .a(N17), .b(N42), .O(N322) );
and2 gate35( .a(N17_OBF), .b(N42), .O(N323) );
nand2 gate36( .a(N159), .b(N165), .O(N324) );
or2 gate37( .a(N159), .b(N165), .O(N325) );
nand2 gate38( .a(N171), .b(N177), .O(N326) );
or2 gate39( .a(N171), .b(N177), .O(N327) );
nand2 gate40( .a(N183), .b(N189), .O(N328) );
or2 gate41( .a(N183), .b(N189), .O(N329) );
nand2 gate42( .a(N195), .b(N201), .O(N330) );
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
and2 gate45( .a(N210), .b(N96), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
and2 gate48( .a(N210), .b(N111), .O(N336) );
and2 gate49( .a(N255), .b(N259), .O(N337) );
and2 gate50( .a(N210), .b(N116), .O(N338) );
and2 gate51( .a(N255_OBF), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
and2 gate53( .a(N255), .b(N267), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
or2 gate56( .a(N270), .b(N273), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );
nor2 gate60( .a(N280), .b(N284), .O(N348) );
or2 gate61( .a(N280), .b(N285), .O(N349) );
or2 gate62( .a(N280), .b(N286), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );
nand2 gate67( .a(N89), .b(N298), .O(N355) );
and2 gate68( .a(N90), .b(N298), .O(N356) );
nand2 gate69( .a(N301), .b(N302), .O(N357) );
nand2 gate70( .a(N303), .b(N304), .O(N360) );
nand2 gate71( .a(N305), .b(N306), .O(N363) );
nand2 gate72( .a(N307), .b(N308), .O(N366) );
inv1 gate73( .a(N310), .O(N369) );
nor2 gate74( .a(N322), .b(N323), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );
nand2 gate76( .a(N326), .b(N327), .O(N379) );
nand2 gate77( .a(N328), .b(N329), .O(N382) );
nand2 gate78( .a(N330), .b(N331), .O(N385) );
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
and2 gate86( .a(N348), .b(N73), .O(N400) );
inv1 gate87( .a(N349_OBF), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
and2 gate92( .a(N357), .b(N360), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
and2 gate95( .a(N363), .b(N366), .O(N409) );
nand2 gate96( .a(N347), .b(N352), .O(N410) );
inv1 gate97( .a(N376_OBF), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
and2 gate103( .a(N210), .b(N369), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
and2 gate112( .a(N407), .b(N408), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
and2 gate118( .a(N411), .b(N412), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );
nor2 gate126( .a(N406), .b(N425), .O(N460) );
nor2 gate127( .a(N409), .b(N426), .O(N463) );
nand2 gate128( .a(N442), .b(N410), .O(N466) );
and2 gate129( .a(N143), .b(N427), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
and2 gate134( .a(N310), .b(N432), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );
nand2 gate137( .a(N443), .b(N1), .O(N483) );
or2 gate138( .a(N369), .b(N437), .O(N488) );
or2 gate139( .a(N369), .b(N437), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );
nor2 gate142( .a(N413), .b(N444), .O(N492) );
nor2 gate143( .a(N416), .b(N445), .O(N495) );
nand2 gate144( .a(N130), .b(N460), .O(N498) );
or2 gate145( .a(N130), .b(N460), .O(N499) );
nand2 gate146( .a(N463), .b(N135), .O(N500) );
or2 gate147( .a(N463), .b(N135), .O(N501) );
and2 gate148( .a(N91), .b(N466), .O(N502) );
nor2 gate149( .a(N475), .b(N476), .O(N503) );
and2 gate150( .a(N96), .b(N466), .O(N504) );
nor2 gate151( .a(N477), .b(N478), .O(N505) );
and2 gate152( .a(N101), .b(N466), .O(N506) );
nor2 gate153( .a(N479), .b(N480), .O(N507) );
and2 gate154( .a(N106), .b(N466), .O(N508) );
nor2 gate155( .a(N481), .b(N482), .O(N509) );
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
and2 gate158( .a(N146), .b(N483), .O(N512) );
and2 gate159( .a(N116), .b(N466), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
and2 gate162( .a(N153), .b(N483), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );
nand2 gate164( .a(N130), .b(N492), .O(N518) );
or2 gate165( .a(N130_OBF), .b(N492), .O(N519) );
nand2 gate166( .a(N495), .b(N207), .O(N520) );
or2 gate167( .a(N495), .b(N207), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
and2 gate169( .a(N451), .b(N165), .O(N523) );
and2 gate170( .a(N451_OBF), .b(N171), .O(N524) );
and2 gate171( .a(N451), .b(N177), .O(N525) );
and2 gate172( .a(N451_OBF), .b(N183), .O(N526) );
nand2 gate173( .a(N451), .b(N189), .O(N527) );
nand2 gate174( .a(N451), .b(N195), .O(N528) );
nand2 gate175( .a(N451), .b(N201), .O(N529) );
nand2 gate176( .a(N498), .b(N499), .O(N530) );
nand2 gate177( .a(N500), .b(N501), .O(N533) );
nor2 gate178( .a(N309), .b(N502), .O(N536) );
nor2 gate179( .a(N316), .b(N504), .O(N537) );
nor2 gate180( .a(N317), .b(N506), .O(N538) );
nor2 gate181( .a(N318), .b(N508), .O(N539) );
nor2 gate182( .a(N510), .b(N511), .O(N540) );
nor2 gate183( .a(N512), .b(N513), .O(N541) );
nor2 gate184( .a(N514), .b(N515), .O(N542) );
nor2 gate185( .a(N516), .b(N517), .O(N543) );
nand2 gate186( .a(N518), .b(N519), .O(N544) );
nand2 gate187( .a(N520), .b(N521), .O(N547) );
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533_OBF), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );
nand2 gate191( .a(N536), .b(N503), .O(N553) );
nand2 gate192( .a(N537), .b(N505), .O(N557) );
nand2 gate193( .a(N538), .b(N507), .O(N561) );
nand2 gate194( .a(N539), .b(N509), .O(N565) );
nand2 gate195( .a(N488), .b(N540), .O(N569) );
nand2 gate196( .a(N489), .b(N541), .O(N573) );
nand2 gate197( .a(N490), .b(N542), .O(N577) );
nand2 gate198( .a(N491), .b(N543), .O(N581) );
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
and2 gate202( .a(N550), .b(N551), .O(N588) );
and2 gate203( .a(N585), .b(N586), .O(N589) );
nand2 gate204( .a(N553), .b(N159), .O(N590) );
or2 gate205( .a(N553), .b(N159), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );
nand2 gate207( .a(N557_OBF), .b(N165), .O(N597) );
or2 gate208( .a(N557), .b(N165), .O(N600) );
and2 gate209( .a(N246), .b(N557), .O(N605) );
nand2 gate210( .a(N561), .b(N171), .O(N606) );
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );
nand2 gate213( .a(N565), .b(N177), .O(N616) );
or2 gate214( .a(N565), .b(N177), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );
nand2 gate216( .a(N569), .b(N183), .O(N625) );
or2 gate217( .a(N569), .b(N183), .O(N628) );
and2 gate218( .a(N246), .b(N569), .O(N631) );
nand2 gate219( .a(N573), .b(N189), .O(N632) );
or2 gate220( .a(N573), .b(N189), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );
nand2 gate222( .a(N577), .b(N195), .O(N641) );
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );
nand2 gate225( .a(N581), .b(N201), .O(N651) );
or2 gate226( .a(N581), .b(N201), .O(N654) );
and2 gate227( .a(N246), .b(N581), .O(N659) );
nor2 gate228( .a(N552), .b(N588), .O(N660) );
nor2 gate229( .a(N587), .b(N589), .O(N661) );
inv1 gate230( .a(N590), .O(N662) );
and2 gate231( .a(N593), .b(N590), .O(N665) );
nor2 gate232( .a(N596), .b(N522), .O(N669) );
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );
nor2 gate235( .a(N605), .b(N523), .O(N677) );
inv1 gate236( .a(N606), .O(N678) );
and2 gate237( .a(N609), .b(N606), .O(N682) );
nor2 gate238( .a(N615), .b(N524), .O(N686) );
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );
nor2 gate241( .a(N624), .b(N525), .O(N696) );
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );
nor2 gate244( .a(N631), .b(N526), .O(N704) );
inv1 gate245( .a(N632), .O(N705) );
and2 gate246( .a(N635), .b(N632), .O(N708) );
nor2 gate247( .a(N337), .b(N640), .O(N712) );
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644_OBF), .b(N641), .O(N717) );
nor2 gate250( .a(N339), .b(N650), .O(N721) );
inv1 gate251( .a(N651), .O(N722) );
and2 gate252( .a(N654), .b(N651), .O(N727) );
nor2 gate253( .a(N341), .b(N659), .O(N731) );
nand2 gate254( .a(N654), .b(N261), .O(N732) );
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
and2 gate258( .a(N228), .b(N665), .O(N736) );
and2 gate259( .a(N237), .b(N662), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
and2 gate264( .a(N228), .b(N682), .O(N742) );
and2 gate265( .a(N237), .b(N678), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
and2 gate268( .a(N237), .b(N687), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
and2 gate270( .a(N228), .b(N700), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
and2 gate273( .a(N228), .b(N708), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228_OBF), .b(N717), .O(N754) );
and2 gate277( .a(N237), .b(N713), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );
nor2 gate279( .a(N727), .b(N261), .O(N757) );
and2 gate280( .a(N727), .b(N261), .O(N758) );
and2 gate281( .a(N228), .b(N727), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );
nand2 gate283( .a(N644), .b(N722), .O(N761) );
nand2 gate284( .a(N635), .b(N713), .O(N762) );
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );
nand2 gate286( .a(N609), .b(N687), .O(N764) );
nand2 gate287( .a(N600), .b(N678), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );
nor2 gate291( .a(N736_OBF), .b(N737), .O(N769) );
nor2 gate292( .a(N739_OBF), .b(N740), .O(N770) );
nor2 gate293( .a(N742), .b(N743), .O(N771) );
nor2 gate294( .a(N745), .b(N746), .O(N772) );
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );
nor2 gate296( .a(N748), .b(N749), .O(N777) );
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );
nor2 gate298( .a(N751), .b(N752), .O(N781) );
nand2 gate299( .a(N756), .b(N732), .O(N782) );
nor2 gate300( .a(N754), .b(N755), .O(N785) );
nor2 gate301( .a(N757), .b(N758), .O(N786) );
nor2 gate302( .a(N759_OBF), .b(N760), .O(N787) );
nor2 gate303( .a(N700), .b(N773), .O(N788) );
and2 gate304( .a(N700), .b(N773), .O(N789) );
nor2 gate305( .a(N708), .b(N778), .O(N790) );
and2 gate306( .a(N708), .b(N778), .O(N791) );
nor2 gate307( .a(N717), .b(N782), .O(N792) );
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );
nand2 gate310( .a(N628), .b(N773), .O(N795) );
nand2 gate311( .a(N795), .b(N747), .O(N796) );
nor2 gate312( .a(N788), .b(N789), .O(N802) );
nor2 gate313( .a(N790), .b(N791), .O(N803) );
nor2 gate314( .a(N792), .b(N793), .O(N804) );
nor2 gate315( .a(N340), .b(N794), .O(N805) );
nor2 gate316( .a(N692), .b(N796), .O(N806) );
and2 gate317( .a(N692), .b(N796), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219_OBF), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );
nand2 gate322( .a(N619), .b(N796), .O(N812) );
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600_OBF), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );
nand2 gate327( .a(N744), .b(N812), .O(N822) );
nor2 gate328( .a(N806), .b(N807), .O(N825) );
nor2 gate329( .a(N335), .b(N808), .O(N826) );
nor2 gate330( .a(N336), .b(N809), .O(N827) );
nor2 gate331( .a(N338), .b(N810), .O(N828) );
inv1 gate332( .a(N811), .O(N829) );
nor2 gate333( .a(N665), .b(N815), .O(N830) );
and2 gate334( .a(N665), .b(N815), .O(N831) );
nor2 gate335( .a(N673), .b(N819), .O(N832) );
and2 gate336( .a(N673), .b(N819), .O(N833) );
nor2 gate337( .a(N682), .b(N822), .O(N834) );
and2 gate338( .a(N682), .b(N822), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );
nand2 gate344( .a(N815), .b(N593), .O(N841) );
nor2 gate345( .a(N830_OBF), .b(N831), .O(N842) );
nor2 gate346( .a(N832), .b(N833), .O(N843) );
nor2 gate347( .a(N834), .b(N835), .O(N844) );
nor2 gate348( .a(N334), .b(N836), .O(N845) );
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
and2 gate354( .a(N219), .b(N842), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );
nor2 gate362( .a(N417_OBF), .b(N851), .O(N859) );
nor2 gate363( .a(N332), .b(N852), .O(N860) );
nor2 gate364( .a(N333), .b(N853), .O(N861) );
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );
inv1 gate( .a(D_0), .O(D_0_NOT) );
inv1 gate( .a(D_1), .O(D_1_NOT) );
inv1 gate( .a(N255), .O(N255_NOT) );
and2 gate( .a(N255), .b(D_0_NOT), .O(ED_0) );
and2 gate( .a(N255_NOT), .b(D_0_NOT), .O(ED_1) );
and2 gate( .a(CONST1), .b(D_0), .O(ED_2) );
and2 gate( .a(CONST0), .b(D_0), .O(ED_3) );
and2 gate( .a(ED_0), .b(D_1_NOT), .O(ED_9) );
and2 gate( .a(ED_1), .b(D_1), .O(ED_7) );
and2 gate( .a(ED_2), .b(D_1_NOT), .O(ED_5) );
and2 gate( .a(ED_3), .b(D_1), .O(ED_4) );
or2  gate( .a(ED_4), .b(ED_5), .O(ED_6) );
or2  gate( .a(ED_6), .b(ED_7), .O(ED_8) );
or2  gate( .a(ED_9), .b(ED_8), .O(N255_OBF) );
inv1 gate( .a(D_2), .O(D_2_NOT) );
inv1 gate( .a(D_3), .O(D_3_NOT) );
inv1 gate( .a(N600), .O(N600_NOT) );
and2 gate( .a(N600), .b(D_2_NOT), .O(ED_10) );
and2 gate( .a(N600_NOT), .b(D_2_NOT), .O(ED_11) );
and2 gate( .a(CONST1), .b(D_2), .O(ED_12) );
and2 gate( .a(CONST0), .b(D_2), .O(ED_13) );
and2 gate( .a(ED_10), .b(D_3_NOT), .O(ED_19) );
and2 gate( .a(ED_11), .b(D_3), .O(ED_17) );
and2 gate( .a(ED_12), .b(D_3_NOT), .O(ED_15) );
and2 gate( .a(ED_13), .b(D_3), .O(ED_14) );
or2  gate( .a(ED_14), .b(ED_15), .O(ED_16) );
or2  gate( .a(ED_16), .b(ED_17), .O(ED_18) );
or2  gate( .a(ED_19), .b(ED_18), .O(N600_OBF) );
inv1 gate( .a(D_4), .O(D_4_NOT) );
inv1 gate( .a(D_5), .O(D_5_NOT) );
inv1 gate( .a(N739), .O(N739_NOT) );
and2 gate( .a(N739), .b(D_4_NOT), .O(ED_20) );
and2 gate( .a(N739_NOT), .b(D_4_NOT), .O(ED_21) );
and2 gate( .a(CONST1), .b(D_4), .O(ED_22) );
and2 gate( .a(CONST0), .b(D_4), .O(ED_23) );
and2 gate( .a(ED_20), .b(D_5_NOT), .O(ED_29) );
and2 gate( .a(ED_21), .b(D_5), .O(ED_27) );
and2 gate( .a(ED_22), .b(D_5_NOT), .O(ED_25) );
and2 gate( .a(ED_23), .b(D_5), .O(ED_24) );
or2  gate( .a(ED_24), .b(ED_25), .O(ED_26) );
or2  gate( .a(ED_26), .b(ED_27), .O(ED_28) );
or2  gate( .a(ED_29), .b(ED_28), .O(N739_OBF) );
inv1 gate( .a(D_6), .O(D_6_NOT) );
inv1 gate( .a(D_7), .O(D_7_NOT) );
inv1 gate( .a(N376), .O(N376_NOT) );
and2 gate( .a(N376), .b(D_6_NOT), .O(ED_30) );
and2 gate( .a(N376_NOT), .b(D_6_NOT), .O(ED_31) );
and2 gate( .a(CONST1), .b(D_6), .O(ED_32) );
and2 gate( .a(CONST0), .b(D_6), .O(ED_33) );
and2 gate( .a(ED_30), .b(D_7_NOT), .O(ED_39) );
and2 gate( .a(ED_31), .b(D_7), .O(ED_37) );
and2 gate( .a(ED_32), .b(D_7_NOT), .O(ED_35) );
and2 gate( .a(ED_33), .b(D_7), .O(ED_34) );
or2  gate( .a(ED_34), .b(ED_35), .O(ED_36) );
or2  gate( .a(ED_36), .b(ED_37), .O(ED_38) );
or2  gate( .a(ED_39), .b(ED_38), .O(N376_OBF) );
inv1 gate( .a(D_8), .O(D_8_NOT) );
inv1 gate( .a(D_9), .O(D_9_NOT) );
inv1 gate( .a(N533), .O(N533_NOT) );
and2 gate( .a(N533), .b(D_8_NOT), .O(ED_40) );
and2 gate( .a(N533_NOT), .b(D_8_NOT), .O(ED_41) );
and2 gate( .a(CONST1), .b(D_8), .O(ED_42) );
and2 gate( .a(CONST0), .b(D_8), .O(ED_43) );
and2 gate( .a(ED_40), .b(D_9_NOT), .O(ED_49) );
and2 gate( .a(ED_41), .b(D_9), .O(ED_47) );
and2 gate( .a(ED_42), .b(D_9_NOT), .O(ED_45) );
and2 gate( .a(ED_43), .b(D_9), .O(ED_44) );
or2  gate( .a(ED_44), .b(ED_45), .O(ED_46) );
or2  gate( .a(ED_46), .b(ED_47), .O(ED_48) );
or2  gate( .a(ED_49), .b(ED_48), .O(N533_OBF) );
inv1 gate( .a(D_10), .O(D_10_NOT) );
inv1 gate( .a(D_11), .O(D_11_NOT) );
inv1 gate( .a(N451), .O(N451_NOT) );
and2 gate( .a(N451), .b(D_10_NOT), .O(ED_50) );
and2 gate( .a(N451_NOT), .b(D_10_NOT), .O(ED_51) );
and2 gate( .a(CONST1), .b(D_10), .O(ED_52) );
and2 gate( .a(CONST0), .b(D_10), .O(ED_53) );
and2 gate( .a(ED_50), .b(D_11_NOT), .O(ED_59) );
and2 gate( .a(ED_51), .b(D_11), .O(ED_57) );
and2 gate( .a(ED_52), .b(D_11_NOT), .O(ED_55) );
and2 gate( .a(ED_53), .b(D_11), .O(ED_54) );
or2  gate( .a(ED_54), .b(ED_55), .O(ED_56) );
or2  gate( .a(ED_56), .b(ED_57), .O(ED_58) );
or2  gate( .a(ED_59), .b(ED_58), .O(N451_OBF) );
inv1 gate( .a(D_12), .O(D_12_NOT) );
inv1 gate( .a(D_13), .O(D_13_NOT) );
inv1 gate( .a(N644), .O(N644_NOT) );
and2 gate( .a(N644), .b(D_12_NOT), .O(ED_60) );
and2 gate( .a(N644_NOT), .b(D_12_NOT), .O(ED_61) );
and2 gate( .a(CONST1), .b(D_12), .O(ED_62) );
and2 gate( .a(CONST0), .b(D_12), .O(ED_63) );
and2 gate( .a(ED_60), .b(D_13_NOT), .O(ED_69) );
and2 gate( .a(ED_61), .b(D_13), .O(ED_67) );
and2 gate( .a(ED_62), .b(D_13_NOT), .O(ED_65) );
and2 gate( .a(ED_63), .b(D_13), .O(ED_64) );
or2  gate( .a(ED_64), .b(ED_65), .O(ED_66) );
or2  gate( .a(ED_66), .b(ED_67), .O(ED_68) );
or2  gate( .a(ED_69), .b(ED_68), .O(N644_OBF) );
inv1 gate( .a(D_14), .O(D_14_NOT) );
inv1 gate( .a(D_15), .O(D_15_NOT) );
inv1 gate( .a(N759), .O(N759_NOT) );
and2 gate( .a(N759), .b(D_14_NOT), .O(ED_70) );
and2 gate( .a(N759_NOT), .b(D_14_NOT), .O(ED_71) );
and2 gate( .a(CONST1), .b(D_14), .O(ED_72) );
and2 gate( .a(CONST0), .b(D_14), .O(ED_73) );
and2 gate( .a(ED_70), .b(D_15_NOT), .O(ED_79) );
and2 gate( .a(ED_71), .b(D_15), .O(ED_77) );
and2 gate( .a(ED_72), .b(D_15_NOT), .O(ED_75) );
and2 gate( .a(ED_73), .b(D_15), .O(ED_74) );
or2  gate( .a(ED_74), .b(ED_75), .O(ED_76) );
or2  gate( .a(ED_76), .b(ED_77), .O(ED_78) );
or2  gate( .a(ED_79), .b(ED_78), .O(N759_OBF) );
inv1 gate( .a(D_16), .O(D_16_NOT) );
inv1 gate( .a(D_17), .O(D_17_NOT) );
inv1 gate( .a(N17), .O(N17_NOT) );
and2 gate( .a(N17), .b(D_16_NOT), .O(ED_80) );
and2 gate( .a(N17_NOT), .b(D_16_NOT), .O(ED_81) );
and2 gate( .a(CONST1), .b(D_16), .O(ED_82) );
and2 gate( .a(CONST0), .b(D_16), .O(ED_83) );
and2 gate( .a(ED_80), .b(D_17_NOT), .O(ED_89) );
and2 gate( .a(ED_81), .b(D_17), .O(ED_87) );
and2 gate( .a(ED_82), .b(D_17_NOT), .O(ED_85) );
and2 gate( .a(ED_83), .b(D_17), .O(ED_84) );
or2  gate( .a(ED_84), .b(ED_85), .O(ED_86) );
or2  gate( .a(ED_86), .b(ED_87), .O(ED_88) );
or2  gate( .a(ED_89), .b(ED_88), .O(N17_OBF) );
inv1 gate( .a(D_18), .O(D_18_NOT) );
inv1 gate( .a(D_19), .O(D_19_NOT) );
inv1 gate( .a(N29), .O(N29_NOT) );
and2 gate( .a(N29), .b(D_18_NOT), .O(ED_90) );
and2 gate( .a(N29_NOT), .b(D_18_NOT), .O(ED_91) );
and2 gate( .a(CONST1), .b(D_18), .O(ED_92) );
and2 gate( .a(CONST0), .b(D_18), .O(ED_93) );
and2 gate( .a(ED_90), .b(D_19_NOT), .O(ED_99) );
and2 gate( .a(ED_91), .b(D_19), .O(ED_97) );
and2 gate( .a(ED_92), .b(D_19_NOT), .O(ED_95) );
and2 gate( .a(ED_93), .b(D_19), .O(ED_94) );
or2  gate( .a(ED_94), .b(ED_95), .O(ED_96) );
or2  gate( .a(ED_96), .b(ED_97), .O(ED_98) );
or2  gate( .a(ED_99), .b(ED_98), .O(N29_OBF) );
inv1 gate( .a(D_20), .O(D_20_NOT) );
inv1 gate( .a(D_21), .O(D_21_NOT) );
inv1 gate( .a(N219), .O(N219_NOT) );
and2 gate( .a(N219), .b(D_20_NOT), .O(ED_100) );
and2 gate( .a(N219_NOT), .b(D_20_NOT), .O(ED_101) );
and2 gate( .a(CONST1), .b(D_20), .O(ED_102) );
and2 gate( .a(CONST0), .b(D_20), .O(ED_103) );
and2 gate( .a(ED_100), .b(D_21_NOT), .O(ED_109) );
and2 gate( .a(ED_101), .b(D_21), .O(ED_107) );
and2 gate( .a(ED_102), .b(D_21_NOT), .O(ED_105) );
and2 gate( .a(ED_103), .b(D_21), .O(ED_104) );
or2  gate( .a(ED_104), .b(ED_105), .O(ED_106) );
or2  gate( .a(ED_106), .b(ED_107), .O(ED_108) );
or2  gate( .a(ED_109), .b(ED_108), .O(N219_OBF) );
inv1 gate( .a(D_22), .O(D_22_NOT) );
inv1 gate( .a(D_23), .O(D_23_NOT) );
inv1 gate( .a(N130), .O(N130_NOT) );
and2 gate( .a(N130), .b(D_22_NOT), .O(ED_110) );
and2 gate( .a(N130_NOT), .b(D_22_NOT), .O(ED_111) );
and2 gate( .a(CONST1), .b(D_22), .O(ED_112) );
and2 gate( .a(CONST0), .b(D_22), .O(ED_113) );
and2 gate( .a(ED_110), .b(D_23_NOT), .O(ED_119) );
and2 gate( .a(ED_111), .b(D_23), .O(ED_117) );
and2 gate( .a(ED_112), .b(D_23_NOT), .O(ED_115) );
and2 gate( .a(ED_113), .b(D_23), .O(ED_114) );
or2  gate( .a(ED_114), .b(ED_115), .O(ED_116) );
or2  gate( .a(ED_116), .b(ED_117), .O(ED_118) );
or2  gate( .a(ED_119), .b(ED_118), .O(N130_OBF) );
inv1 gate( .a(D_24), .O(D_24_NOT) );
inv1 gate( .a(D_25), .O(D_25_NOT) );
inv1 gate( .a(N736), .O(N736_NOT) );
and2 gate( .a(N736), .b(D_24_NOT), .O(ED_120) );
and2 gate( .a(N736_NOT), .b(D_24_NOT), .O(ED_121) );
and2 gate( .a(CONST1), .b(D_24), .O(ED_122) );
and2 gate( .a(CONST0), .b(D_24), .O(ED_123) );
and2 gate( .a(ED_120), .b(D_25_NOT), .O(ED_129) );
and2 gate( .a(ED_121), .b(D_25), .O(ED_127) );
and2 gate( .a(ED_122), .b(D_25_NOT), .O(ED_125) );
and2 gate( .a(ED_123), .b(D_25), .O(ED_124) );
or2  gate( .a(ED_124), .b(ED_125), .O(ED_126) );
or2  gate( .a(ED_126), .b(ED_127), .O(ED_128) );
or2  gate( .a(ED_129), .b(ED_128), .O(N736_OBF) );
inv1 gate( .a(D_26), .O(D_26_NOT) );
inv1 gate( .a(D_27), .O(D_27_NOT) );
inv1 gate( .a(N451), .O(N451_NOT) );
and2 gate( .a(N451), .b(D_26_NOT), .O(ED_130) );
and2 gate( .a(N451_NOT), .b(D_26_NOT), .O(ED_131) );
and2 gate( .a(CONST1), .b(D_26), .O(ED_132) );
and2 gate( .a(CONST0), .b(D_26), .O(ED_133) );
and2 gate( .a(ED_130), .b(D_27_NOT), .O(ED_139) );
and2 gate( .a(ED_131), .b(D_27), .O(ED_137) );
and2 gate( .a(ED_132), .b(D_27_NOT), .O(ED_135) );
and2 gate( .a(ED_133), .b(D_27), .O(ED_134) );
or2  gate( .a(ED_134), .b(ED_135), .O(ED_136) );
or2  gate( .a(ED_136), .b(ED_137), .O(ED_138) );
or2  gate( .a(ED_139), .b(ED_138), .O(N451_OBF) );
inv1 gate( .a(D_28), .O(D_28_NOT) );
inv1 gate( .a(D_29), .O(D_29_NOT) );
inv1 gate( .a(N228), .O(N228_NOT) );
and2 gate( .a(N228), .b(D_28_NOT), .O(ED_140) );
and2 gate( .a(N228_NOT), .b(D_28_NOT), .O(ED_141) );
and2 gate( .a(CONST1), .b(D_28), .O(ED_142) );
and2 gate( .a(CONST0), .b(D_28), .O(ED_143) );
and2 gate( .a(ED_140), .b(D_29_NOT), .O(ED_149) );
and2 gate( .a(ED_141), .b(D_29), .O(ED_147) );
and2 gate( .a(ED_142), .b(D_29_NOT), .O(ED_145) );
and2 gate( .a(ED_143), .b(D_29), .O(ED_144) );
or2  gate( .a(ED_144), .b(ED_145), .O(ED_146) );
or2  gate( .a(ED_146), .b(ED_147), .O(ED_148) );
or2  gate( .a(ED_149), .b(ED_148), .O(N228_OBF) );
inv1 gate( .a(D_30), .O(D_30_NOT) );
inv1 gate( .a(D_31), .O(D_31_NOT) );
inv1 gate( .a(N349), .O(N349_NOT) );
and2 gate( .a(N349), .b(D_30_NOT), .O(ED_150) );
and2 gate( .a(N349_NOT), .b(D_30_NOT), .O(ED_151) );
and2 gate( .a(CONST1), .b(D_30), .O(ED_152) );
and2 gate( .a(CONST0), .b(D_30), .O(ED_153) );
and2 gate( .a(ED_150), .b(D_31_NOT), .O(ED_159) );
and2 gate( .a(ED_151), .b(D_31), .O(ED_157) );
and2 gate( .a(ED_152), .b(D_31_NOT), .O(ED_155) );
and2 gate( .a(ED_153), .b(D_31), .O(ED_154) );
or2  gate( .a(ED_154), .b(ED_155), .O(ED_156) );
or2  gate( .a(ED_156), .b(ED_157), .O(ED_158) );
or2  gate( .a(ED_159), .b(ED_158), .O(N349_OBF) );
inv1 gate( .a(D_32), .O(D_32_NOT) );
inv1 gate( .a(D_33), .O(D_33_NOT) );
inv1 gate( .a(N417), .O(N417_NOT) );
and2 gate( .a(N417), .b(D_32_NOT), .O(ED_160) );
and2 gate( .a(N417_NOT), .b(D_32_NOT), .O(ED_161) );
and2 gate( .a(CONST1), .b(D_32), .O(ED_162) );
and2 gate( .a(CONST0), .b(D_32), .O(ED_163) );
and2 gate( .a(ED_160), .b(D_33_NOT), .O(ED_169) );
and2 gate( .a(ED_161), .b(D_33), .O(ED_167) );
and2 gate( .a(ED_162), .b(D_33_NOT), .O(ED_165) );
and2 gate( .a(ED_163), .b(D_33), .O(ED_164) );
or2  gate( .a(ED_164), .b(ED_165), .O(ED_166) );
or2  gate( .a(ED_166), .b(ED_167), .O(ED_168) );
or2  gate( .a(ED_169), .b(ED_168), .O(N417_OBF) );
inv1 gate( .a(D_34), .O(D_34_NOT) );
inv1 gate( .a(D_35), .O(D_35_NOT) );
inv1 gate( .a(N830), .O(N830_NOT) );
and2 gate( .a(N830), .b(D_34_NOT), .O(ED_170) );
and2 gate( .a(N830_NOT), .b(D_34_NOT), .O(ED_171) );
and2 gate( .a(CONST1), .b(D_34), .O(ED_172) );
and2 gate( .a(CONST0), .b(D_34), .O(ED_173) );
and2 gate( .a(ED_170), .b(D_35_NOT), .O(ED_179) );
and2 gate( .a(ED_171), .b(D_35), .O(ED_177) );
and2 gate( .a(ED_172), .b(D_35_NOT), .O(ED_175) );
and2 gate( .a(ED_173), .b(D_35), .O(ED_174) );
or2  gate( .a(ED_174), .b(ED_175), .O(ED_176) );
or2  gate( .a(ED_176), .b(ED_177), .O(ED_178) );
or2  gate( .a(ED_179), .b(ED_178), .O(N830_OBF) );
inv1 gate( .a(D_36), .O(D_36_NOT) );
inv1 gate( .a(D_37), .O(D_37_NOT) );
inv1 gate( .a(N29), .O(N29_NOT) );
and2 gate( .a(N29), .b(D_36_NOT), .O(ED_180) );
and2 gate( .a(N29_NOT), .b(D_36_NOT), .O(ED_181) );
and2 gate( .a(CONST1), .b(D_36), .O(ED_182) );
and2 gate( .a(CONST0), .b(D_36), .O(ED_183) );
and2 gate( .a(ED_180), .b(D_37_NOT), .O(ED_189) );
and2 gate( .a(ED_181), .b(D_37), .O(ED_187) );
and2 gate( .a(ED_182), .b(D_37_NOT), .O(ED_185) );
and2 gate( .a(ED_183), .b(D_37), .O(ED_184) );
or2  gate( .a(ED_184), .b(ED_185), .O(ED_186) );
or2  gate( .a(ED_186), .b(ED_187), .O(ED_188) );
or2  gate( .a(ED_189), .b(ED_188), .O(N29_OBF) );
inv1 gate( .a(D_38), .O(D_38_NOT) );
inv1 gate( .a(D_39), .O(D_39_NOT) );
inv1 gate( .a(N59), .O(N59_NOT) );
and2 gate( .a(N59), .b(D_38_NOT), .O(ED_190) );
and2 gate( .a(N59_NOT), .b(D_38_NOT), .O(ED_191) );
and2 gate( .a(CONST1), .b(D_38), .O(ED_192) );
and2 gate( .a(CONST0), .b(D_38), .O(ED_193) );
and2 gate( .a(ED_190), .b(D_39_NOT), .O(ED_199) );
and2 gate( .a(ED_191), .b(D_39), .O(ED_197) );
and2 gate( .a(ED_192), .b(D_39_NOT), .O(ED_195) );
and2 gate( .a(ED_193), .b(D_39), .O(ED_194) );
or2  gate( .a(ED_194), .b(ED_195), .O(ED_196) );
or2  gate( .a(ED_196), .b(ED_197), .O(ED_198) );
or2  gate( .a(ED_199), .b(ED_198), .O(N59_OBF) );
inv1 gate( .a(D_40), .O(D_40_NOT) );
inv1 gate( .a(D_41), .O(D_41_NOT) );
inv1 gate( .a(N557), .O(N557_NOT) );
and2 gate( .a(N557), .b(D_40_NOT), .O(ED_200) );
and2 gate( .a(N557_NOT), .b(D_40_NOT), .O(ED_201) );
and2 gate( .a(CONST1), .b(D_40), .O(ED_202) );
and2 gate( .a(CONST0), .b(D_40), .O(ED_203) );
and2 gate( .a(ED_200), .b(D_41_NOT), .O(ED_209) );
and2 gate( .a(ED_201), .b(D_41), .O(ED_207) );
and2 gate( .a(ED_202), .b(D_41_NOT), .O(ED_205) );
and2 gate( .a(ED_203), .b(D_41), .O(ED_204) );
or2  gate( .a(ED_204), .b(ED_205), .O(ED_206) );
or2  gate( .a(ED_206), .b(ED_207), .O(ED_208) );
or2  gate( .a(ED_209), .b(ED_208), .O(N557_OBF) );

endmodule
