module	c17 (N1,N2,N3,N4,N5,N6,N7,N8,N9,N12,N13,N14);

input  N1,N2,N3,N4,N5,CONST1,CONST0 //RE__PI;

input D_0,D_1,D_2,D_3,D_4,D_5,D_6,D_7,D_8,D_9,D_10,D_11,D_12,D_13,D_14,D_15,D_16,D_17,D_18,D_19,D_20,D_21,D_22,D_23,D_24,D_25,D_26,D_27,D_28,D_29 //RE__ALLOW(00,01,10,11);
 
output N10,N11;

wire N6,N7,N8,N9,D_0_NOT,D_1_NOT,N1_NOT,N1_OBF,ED_0,ED_1,ED_2,ED_3,ED_4,ED_5,ED_6,ED_7,ED_8,ED_9,
D_2_NOT,D_3_NOT,N3_NOT,N3_OBF,ED_9,ED_10,ED_11,ED_12,ED_13,ED_14,ED_15,ED_16,ED_17,ED_18,
D_4_NOT,D_5_NOT,N2_NOT,N2_OBF,ED_18,ED_19,ED_20,ED_21,ED_22,ED_23,ED_24,ED_25,ED_26,ED_27,
D_6_NOT,D_7_NOT,N1_NOT,N1_OBF,ED_27,ED_28,ED_29,ED_30,ED_31,ED_32,ED_33,ED_34,ED_35,ED_36,
D_8_NOT,D_9_NOT,N6_OBF_NOT,N6_OBF,ED_36,ED_37,ED_38,ED_39,ED_40,ED_41,ED_42,ED_43,ED_44,ED_45,
D_10_NOT,D_11_NOT,N7_NOT,N7_OBF,ED_45,ED_46,ED_47,ED_48,ED_49,ED_50,ED_51,ED_52,ED_53,ED_54,
D_12_NOT,D_13_NOT,N9_NOT,N9_OBF,ED_54,ED_55,ED_56,ED_57,ED_58,ED_59,ED_60,ED_61,ED_62,ED_63,
D_14_NOT,D_15_NOT,N2_NOT,N2_OBF,ED_63,ED_64,ED_65,ED_66,ED_67,ED_68,ED_69,ED_70,ED_71,ED_72,
D_16_NOT,D_17_NOT,N1_NOT,N1_OBF,ED_72,ED_73,ED_74,ED_75,ED_76,ED_77,ED_78,ED_79,ED_80,ED_81,
D_18_NOT,D_19_NOT,N11_OBF_NOT,N11_OBF,ED_81,ED_82,ED_83,ED_84,ED_85,ED_86,ED_87,ED_88,ED_89,ED_90,
D_20_NOT,D_21_NOT,N6_NOT,N6_OBF,ED_90,ED_91,ED_92,ED_93,ED_94,ED_95,ED_96,ED_97,ED_98,ED_99,
D_22_NOT,D_23_NOT,N7_NOT,N7_OBF,ED_99,ED_100,ED_101,ED_102,ED_103,ED_104,ED_105,ED_106,ED_107,ED_108,
D_24_NOT,D_25_NOT,N2_NOT,N2_OBF,ED_108,ED_109,ED_110,ED_111,ED_112,ED_113,ED_114,ED_115,ED_116,ED_117,
D_26_NOT,D_27_NOT,N1_NOT,N1_OBF,ED_117,ED_118,ED_119,ED_120,ED_121,ED_122,ED_123,ED_124,ED_125,ED_126,
D_28_NOT,D_29_NOT,N10_OBF_NOT,N10_OBF,ED_126,ED_127,ED_128,ED_129,ED_130,ED_131,ED_132,ED_133,ED_134,ED_135;
     
nand2 gate1( .a(N1), .b(N3), .O(N6) );
nand2 gate2( .a(N3), .b(N4), .O(N8) );
nand2 gate3( .a(N2), .b(N8), .O(N7) );
nand2 gate4( .a(N8), .b(N5), .O(N9) );
;
;
inv1 gate( .a(D_0), .O(D_0_NOT) );
inv1 gate( .a(D_1), .O(D_1_NOT) );
inv1 gate( .a(N1), .O(N1_NOT) );
and2 gate( .a(N1), .b(D_0_NOT), .O(ED_0) );
and2 gate( .a(N1_NOT), .b(D_0_NOT), .O(ED_1) );
and2 gate( .a(CONST1), .b(D_0), .O(ED_2) );
and2 gate( .a(CONST0), .b(D_0), .O(ED_3) );
and2 gate( .a(ED_0), .b(D_1_NOT), .O(ED_9) );
and2 gate( .a(ED_1), .b(D_1), .O(ED_7) );
and2 gate( .a(ED_2), .b(D_1_NOT), .O(ED_5) );
and2 gate( .a(ED_3), .b(D_1), .O(ED_4) );
or2  gate( .a(ED_4), .b(ED_5), .O(ED_6) );
or2  gate( .a(ED_6), .b(ED_7), .O(ED_8) );
or2  gate( .a(ED_9), .b(ED_8), .O(N1_OBF);
inv1 gate( .a(D_2), .O(D_2_NOT) );
inv1 gate( .a(D_3), .O(D_3_NOT) );
inv1 gate( .a(N3), .O(N3_NOT) );
and2 gate( .a(N3), .b(D_2_NOT), .O(ED_9) );
and2 gate( .a(N3_NOT), .b(D_2_NOT), .O(ED_10) );
and2 gate( .a(CONST1), .b(D_2), .O(ED_11) );
and2 gate( .a(CONST0), .b(D_2), .O(ED_12) );
and2 gate( .a(ED_9), .b(D_3_NOT), .O(ED_18) );
and2 gate( .a(ED_10), .b(D_3), .O(ED_16) );
and2 gate( .a(ED_11), .b(D_3_NOT), .O(ED_14) );
and2 gate( .a(ED_12), .b(D_3), .O(ED_13) );
or2  gate( .a(ED_13), .b(ED_14), .O(ED_15) );
or2  gate( .a(ED_15), .b(ED_16), .O(ED_17) );
or2  gate( .a(ED_18), .b(ED_17), .O(N3_OBF);
inv1 gate( .a(D_4), .O(D_4_NOT) );
inv1 gate( .a(D_5), .O(D_5_NOT) );
inv1 gate( .a(N2), .O(N2_NOT) );
and2 gate( .a(N2), .b(D_4_NOT), .O(ED_18) );
and2 gate( .a(N2_NOT), .b(D_4_NOT), .O(ED_19) );
and2 gate( .a(CONST1), .b(D_4), .O(ED_20) );
and2 gate( .a(CONST0), .b(D_4), .O(ED_21) );
and2 gate( .a(ED_18), .b(D_5_NOT), .O(ED_27) );
and2 gate( .a(ED_19), .b(D_5), .O(ED_25) );
and2 gate( .a(ED_20), .b(D_5_NOT), .O(ED_23) );
and2 gate( .a(ED_21), .b(D_5), .O(ED_22) );
or2  gate( .a(ED_22), .b(ED_23), .O(ED_24) );
or2  gate( .a(ED_24), .b(ED_25), .O(ED_26) );
or2  gate( .a(ED_27), .b(ED_26), .O(N2_OBF);
inv1 gate( .a(D_6), .O(D_6_NOT) );
inv1 gate( .a(D_7), .O(D_7_NOT) );
inv1 gate( .a(N1), .O(N1_NOT) );
and2 gate( .a(N1), .b(D_6_NOT), .O(ED_27) );
and2 gate( .a(N1_NOT), .b(D_6_NOT), .O(ED_28) );
and2 gate( .a(CONST1), .b(D_6), .O(ED_29) );
and2 gate( .a(CONST0), .b(D_6), .O(ED_30) );
and2 gate( .a(ED_27), .b(D_7_NOT), .O(ED_36) );
and2 gate( .a(ED_28), .b(D_7), .O(ED_34) );
and2 gate( .a(ED_29), .b(D_7_NOT), .O(ED_32) );
and2 gate( .a(ED_30), .b(D_7), .O(ED_31) );
or2  gate( .a(ED_31), .b(ED_32), .O(ED_33) );
or2  gate( .a(ED_33), .b(ED_34), .O(ED_35) );
or2  gate( .a(ED_36), .b(ED_35), .O(N1_OBF);
inv1 gate( .a(D_8), .O(D_8_NOT) );
inv1 gate( .a(D_9), .O(D_9_NOT) );
inv1 gate( .a(N6_OBF), .O(N6_OBF_NOT) );
and2 gate( .a(N6_OBF), .b(D_8_NOT), .O(ED_36) );
and2 gate( .a(N6_OBF_NOT), .b(D_8_NOT), .O(ED_37) );
and2 gate( .a(CONST1), .b(D_8), .O(ED_38) );
and2 gate( .a(CONST0), .b(D_8), .O(ED_39) );
and2 gate( .a(ED_36), .b(D_9_NOT), .O(ED_45) );
and2 gate( .a(ED_37), .b(D_9), .O(ED_43) );
and2 gate( .a(ED_38), .b(D_9_NOT), .O(ED_41) );
and2 gate( .a(ED_39), .b(D_9), .O(ED_40) );
or2  gate( .a(ED_40), .b(ED_41), .O(ED_42) );
or2  gate( .a(ED_42), .b(ED_43), .O(ED_44) );
or2  gate( .a(ED_45), .b(ED_44), .O(N6);
nand4 gate( .a(N1_OBF), .b(N3_OBF), .c(N2_OBF), .d(N1_OBF), .O(N6_OBF) );
inv1 gate( .a(D_10), .O(D_10_NOT) );
inv1 gate( .a(D_11), .O(D_11_NOT) );
inv1 gate( .a(N7), .O(N7_NOT) );
and2 gate( .a(N7), .b(D_10_NOT), .O(ED_45) );
and2 gate( .a(N7_NOT), .b(D_10_NOT), .O(ED_46) );
and2 gate( .a(CONST1), .b(D_10), .O(ED_47) );
and2 gate( .a(CONST0), .b(D_10), .O(ED_48) );
and2 gate( .a(ED_45), .b(D_11_NOT), .O(ED_54) );
and2 gate( .a(ED_46), .b(D_11), .O(ED_52) );
and2 gate( .a(ED_47), .b(D_11_NOT), .O(ED_50) );
and2 gate( .a(ED_48), .b(D_11), .O(ED_49) );
or2  gate( .a(ED_49), .b(ED_50), .O(ED_51) );
or2  gate( .a(ED_51), .b(ED_52), .O(ED_53) );
or2  gate( .a(ED_54), .b(ED_53), .O(N7_OBF);
inv1 gate( .a(D_12), .O(D_12_NOT) );
inv1 gate( .a(D_13), .O(D_13_NOT) );
inv1 gate( .a(N9), .O(N9_NOT) );
and2 gate( .a(N9), .b(D_12_NOT), .O(ED_54) );
and2 gate( .a(N9_NOT), .b(D_12_NOT), .O(ED_55) );
and2 gate( .a(CONST1), .b(D_12), .O(ED_56) );
and2 gate( .a(CONST0), .b(D_12), .O(ED_57) );
and2 gate( .a(ED_54), .b(D_13_NOT), .O(ED_63) );
and2 gate( .a(ED_55), .b(D_13), .O(ED_61) );
and2 gate( .a(ED_56), .b(D_13_NOT), .O(ED_59) );
and2 gate( .a(ED_57), .b(D_13), .O(ED_58) );
or2  gate( .a(ED_58), .b(ED_59), .O(ED_60) );
or2  gate( .a(ED_60), .b(ED_61), .O(ED_62) );
or2  gate( .a(ED_63), .b(ED_62), .O(N9_OBF);
inv1 gate( .a(D_14), .O(D_14_NOT) );
inv1 gate( .a(D_15), .O(D_15_NOT) );
inv1 gate( .a(N2), .O(N2_NOT) );
and2 gate( .a(N2), .b(D_14_NOT), .O(ED_63) );
and2 gate( .a(N2_NOT), .b(D_14_NOT), .O(ED_64) );
and2 gate( .a(CONST1), .b(D_14), .O(ED_65) );
and2 gate( .a(CONST0), .b(D_14), .O(ED_66) );
and2 gate( .a(ED_63), .b(D_15_NOT), .O(ED_72) );
and2 gate( .a(ED_64), .b(D_15), .O(ED_70) );
and2 gate( .a(ED_65), .b(D_15_NOT), .O(ED_68) );
and2 gate( .a(ED_66), .b(D_15), .O(ED_67) );
or2  gate( .a(ED_67), .b(ED_68), .O(ED_69) );
or2  gate( .a(ED_69), .b(ED_70), .O(ED_71) );
or2  gate( .a(ED_72), .b(ED_71), .O(N2_OBF);
inv1 gate( .a(D_16), .O(D_16_NOT) );
inv1 gate( .a(D_17), .O(D_17_NOT) );
inv1 gate( .a(N1), .O(N1_NOT) );
and2 gate( .a(N1), .b(D_16_NOT), .O(ED_72) );
and2 gate( .a(N1_NOT), .b(D_16_NOT), .O(ED_73) );
and2 gate( .a(CONST1), .b(D_16), .O(ED_74) );
and2 gate( .a(CONST0), .b(D_16), .O(ED_75) );
and2 gate( .a(ED_72), .b(D_17_NOT), .O(ED_81) );
and2 gate( .a(ED_73), .b(D_17), .O(ED_79) );
and2 gate( .a(ED_74), .b(D_17_NOT), .O(ED_77) );
and2 gate( .a(ED_75), .b(D_17), .O(ED_76) );
or2  gate( .a(ED_76), .b(ED_77), .O(ED_78) );
or2  gate( .a(ED_78), .b(ED_79), .O(ED_80) );
or2  gate( .a(ED_81), .b(ED_80), .O(N1_OBF);
inv1 gate( .a(D_18), .O(D_18_NOT) );
inv1 gate( .a(D_19), .O(D_19_NOT) );
inv1 gate( .a(N11_OBF), .O(N11_OBF_NOT) );
and2 gate( .a(N11_OBF), .b(D_18_NOT), .O(ED_81) );
and2 gate( .a(N11_OBF_NOT), .b(D_18_NOT), .O(ED_82) );
and2 gate( .a(CONST1), .b(D_18), .O(ED_83) );
and2 gate( .a(CONST0), .b(D_18), .O(ED_84) );
and2 gate( .a(ED_81), .b(D_19_NOT), .O(ED_90) );
and2 gate( .a(ED_82), .b(D_19), .O(ED_88) );
and2 gate( .a(ED_83), .b(D_19_NOT), .O(ED_86) );
and2 gate( .a(ED_84), .b(D_19), .O(ED_85) );
or2  gate( .a(ED_85), .b(ED_86), .O(ED_87) );
or2  gate( .a(ED_87), .b(ED_88), .O(ED_89) );
or2  gate( .a(ED_90), .b(ED_89), .O(N11);
nand4 gate( .a(N7_OBF), .b(N9_OBF), .c(N2_OBF), .d(N1_OBF), .O(N11_OBF) );
inv1 gate( .a(D_20), .O(D_20_NOT) );
inv1 gate( .a(D_21), .O(D_21_NOT) );
inv1 gate( .a(N6), .O(N6_NOT) );
and2 gate( .a(N6), .b(D_20_NOT), .O(ED_90) );
and2 gate( .a(N6_NOT), .b(D_20_NOT), .O(ED_91) );
and2 gate( .a(CONST1), .b(D_20), .O(ED_92) );
and2 gate( .a(CONST0), .b(D_20), .O(ED_93) );
and2 gate( .a(ED_90), .b(D_21_NOT), .O(ED_99) );
and2 gate( .a(ED_91), .b(D_21), .O(ED_97) );
and2 gate( .a(ED_92), .b(D_21_NOT), .O(ED_95) );
and2 gate( .a(ED_93), .b(D_21), .O(ED_94) );
or2  gate( .a(ED_94), .b(ED_95), .O(ED_96) );
or2  gate( .a(ED_96), .b(ED_97), .O(ED_98) );
or2  gate( .a(ED_99), .b(ED_98), .O(N6_OBF);
inv1 gate( .a(D_22), .O(D_22_NOT) );
inv1 gate( .a(D_23), .O(D_23_NOT) );
inv1 gate( .a(N7), .O(N7_NOT) );
and2 gate( .a(N7), .b(D_22_NOT), .O(ED_99) );
and2 gate( .a(N7_NOT), .b(D_22_NOT), .O(ED_100) );
and2 gate( .a(CONST1), .b(D_22), .O(ED_101) );
and2 gate( .a(CONST0), .b(D_22), .O(ED_102) );
and2 gate( .a(ED_99), .b(D_23_NOT), .O(ED_108) );
and2 gate( .a(ED_100), .b(D_23), .O(ED_106) );
and2 gate( .a(ED_101), .b(D_23_NOT), .O(ED_104) );
and2 gate( .a(ED_102), .b(D_23), .O(ED_103) );
or2  gate( .a(ED_103), .b(ED_104), .O(ED_105) );
or2  gate( .a(ED_105), .b(ED_106), .O(ED_107) );
or2  gate( .a(ED_108), .b(ED_107), .O(N7_OBF);
inv1 gate( .a(D_24), .O(D_24_NOT) );
inv1 gate( .a(D_25), .O(D_25_NOT) );
inv1 gate( .a(N2), .O(N2_NOT) );
and2 gate( .a(N2), .b(D_24_NOT), .O(ED_108) );
and2 gate( .a(N2_NOT), .b(D_24_NOT), .O(ED_109) );
and2 gate( .a(CONST1), .b(D_24), .O(ED_110) );
and2 gate( .a(CONST0), .b(D_24), .O(ED_111) );
and2 gate( .a(ED_108), .b(D_25_NOT), .O(ED_117) );
and2 gate( .a(ED_109), .b(D_25), .O(ED_115) );
and2 gate( .a(ED_110), .b(D_25_NOT), .O(ED_113) );
and2 gate( .a(ED_111), .b(D_25), .O(ED_112) );
or2  gate( .a(ED_112), .b(ED_113), .O(ED_114) );
or2  gate( .a(ED_114), .b(ED_115), .O(ED_116) );
or2  gate( .a(ED_117), .b(ED_116), .O(N2_OBF);
inv1 gate( .a(D_26), .O(D_26_NOT) );
inv1 gate( .a(D_27), .O(D_27_NOT) );
inv1 gate( .a(N1), .O(N1_NOT) );
and2 gate( .a(N1), .b(D_26_NOT), .O(ED_117) );
and2 gate( .a(N1_NOT), .b(D_26_NOT), .O(ED_118) );
and2 gate( .a(CONST1), .b(D_26), .O(ED_119) );
and2 gate( .a(CONST0), .b(D_26), .O(ED_120) );
and2 gate( .a(ED_117), .b(D_27_NOT), .O(ED_126) );
and2 gate( .a(ED_118), .b(D_27), .O(ED_124) );
and2 gate( .a(ED_119), .b(D_27_NOT), .O(ED_122) );
and2 gate( .a(ED_120), .b(D_27), .O(ED_121) );
or2  gate( .a(ED_121), .b(ED_122), .O(ED_123) );
or2  gate( .a(ED_123), .b(ED_124), .O(ED_125) );
or2  gate( .a(ED_126), .b(ED_125), .O(N1_OBF);
inv1 gate( .a(D_28), .O(D_28_NOT) );
inv1 gate( .a(D_29), .O(D_29_NOT) );
inv1 gate( .a(N10_OBF), .O(N10_OBF_NOT) );
and2 gate( .a(N10_OBF), .b(D_28_NOT), .O(ED_126) );
and2 gate( .a(N10_OBF_NOT), .b(D_28_NOT), .O(ED_127) );
and2 gate( .a(CONST1), .b(D_28), .O(ED_128) );
and2 gate( .a(CONST0), .b(D_28), .O(ED_129) );
and2 gate( .a(ED_126), .b(D_29_NOT), .O(ED_135) );
and2 gate( .a(ED_127), .b(D_29), .O(ED_133) );
and2 gate( .a(ED_128), .b(D_29_NOT), .O(ED_131) );
and2 gate( .a(ED_129), .b(D_29), .O(ED_130) );
or2  gate( .a(ED_130), .b(ED_131), .O(ED_132) );
or2  gate( .a(ED_132), .b(ED_133), .O(ED_134) );
or2  gate( .a(ED_135), .b(ED_134), .O(N10);
nand4 gate( .a(N6_OBF), .b(N7_OBF), .c(N2_OBF), .d(N1_OBF), .O(N10_OBF) );

endmodule
