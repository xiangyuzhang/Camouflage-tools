
module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input  N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,      N99,N102,N105,N108,N112,N115,CONST1,CONST0 //RE__PI;

input D_0,D_1,D_2,D_3,D_4,D_5,D_6,D_7,D_8,D_9,D_10,D_11,D_12,D_13,D_14,D_15,D_16,D_17,D_18,D_19 //RE__ALLOW(00,01,10,11);

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429,D_0_NOT,D_1_NOT,N246_NOT,N246_OBF,ED_0,ED_1,ED_2,ED_3,ED_4,ED_5,ED_6,ED_7,ED_8,ED_9,D_2_NOT,D_3_NOT,N336_NOT,N336_OBF,ED_9,ED_10,ED_11,ED_12,ED_13,ED_14,ED_15,ED_16,ED_17,ED_18,D_4_NOT,D_5_NOT,N372_NOT,N372_OBF,ED_18,ED_19,ED_20,ED_21,ED_22,ED_23,ED_24,ED_25,ED_26,ED_27,D_6_NOT,D_7_NOT,N17_NOT,N17_OBF,ED_27,ED_28,ED_29,ED_30,ED_31,ED_32,ED_33,ED_34,ED_35,ED_36,D_8_NOT,D_9_NOT,N381_NOT,N381_OBF,ED_36,ED_37,ED_38,ED_39,ED_40,ED_41,ED_42,ED_43,ED_44,ED_45,D_10_NOT,D_11_NOT,N381_NOT,N381_OBF,ED_45,ED_46,ED_47,ED_48,ED_49,ED_50,ED_51,ED_52,ED_53,ED_54,D_12_NOT,D_13_NOT,N386_NOT,N386_OBF,ED_54,ED_55,ED_56,ED_57,ED_58,ED_59,ED_60,ED_61,ED_62,ED_63,D_14_NOT,D_15_NOT,N422_NOT,N422_OBF,ED_63,ED_64,ED_65,ED_66,ED_67,ED_68,ED_69,ED_70,ED_71,ED_72,D_16_NOT,D_17_NOT,N399_NOT,N399_OBF,ED_72,ED_73,ED_74,ED_75,ED_76,ED_77,ED_78,ED_79,ED_80,ED_81,D_18_NOT,D_19_NOT,N430_NOT,N430_OBF,ED_81,ED_82,ED_83,ED_84,ED_85,ED_86,ED_87,ED_88,ED_89,ED_90;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246_OBF), .b(N336_OBF), .c(N372_OBF), .d(N17_OBF), .O(N381_OBF) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381_OBF), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381_OBF), .b(N386), .c(N422), .d(N399), .O(N430_OBF) );
nand4 gate159( .a(N381_OBF), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381_OBF), .b(N422), .c(N425), .d(N429), .O(N432) );
inv1 gate( .a(D_0), .O(D_0_NOT) );
inv1 gate( .a(D_1), .O(D_1_NOT) );
inv1 gate( .a(N246), .O(N246_NOT) );
and2 gate( .a(N246), .b(D_0_NOT), .O(ED_0) );
and2 gate( .a(N246_NOT), .b(D_0_NOT), .O(ED_1) );
and2 gate( .a(CONST1), .b(D_0), .O(ED_2) );
and2 gate( .a(CONST0), .b(D_0), .O(ED_3) );
and2 gate( .a(ED_0), .b(D_1_NOT), .O(ED_9) );
and2 gate( .a(ED_1), .b(D_1), .O(ED_7) );
and2 gate( .a(ED_2), .b(D_1_NOT), .O(ED_5) );
and2 gate( .a(ED_3), .b(D_1), .O(ED_4) );
or2  gate( .a(ED_4), .b(ED_5), .O(ED_6) );
or2  gate( .a(ED_6), .b(ED_7), .O(ED_8) );
or2  gate( .a(ED_9), .b(ED_8), .O(N246_OBF);
inv1 gate( .a(D_2), .O(D_2_NOT) );
inv1 gate( .a(D_3), .O(D_3_NOT) );
inv1 gate( .a(N336), .O(N336_NOT) );
and2 gate( .a(N336), .b(D_2_NOT), .O(ED_9) );
and2 gate( .a(N336_NOT), .b(D_2_NOT), .O(ED_10) );
and2 gate( .a(CONST1), .b(D_2), .O(ED_11) );
and2 gate( .a(CONST0), .b(D_2), .O(ED_12) );
and2 gate( .a(ED_9), .b(D_3_NOT), .O(ED_18) );
and2 gate( .a(ED_10), .b(D_3), .O(ED_16) );
and2 gate( .a(ED_11), .b(D_3_NOT), .O(ED_14) );
and2 gate( .a(ED_12), .b(D_3), .O(ED_13) );
or2  gate( .a(ED_13), .b(ED_14), .O(ED_15) );
or2  gate( .a(ED_15), .b(ED_16), .O(ED_17) );
or2  gate( .a(ED_18), .b(ED_17), .O(N336_OBF);
inv1 gate( .a(D_4), .O(D_4_NOT) );
inv1 gate( .a(D_5), .O(D_5_NOT) );
inv1 gate( .a(N372), .O(N372_NOT) );
and2 gate( .a(N372), .b(D_4_NOT), .O(ED_18) );
and2 gate( .a(N372_NOT), .b(D_4_NOT), .O(ED_19) );
and2 gate( .a(CONST1), .b(D_4), .O(ED_20) );
and2 gate( .a(CONST0), .b(D_4), .O(ED_21) );
and2 gate( .a(ED_18), .b(D_5_NOT), .O(ED_27) );
and2 gate( .a(ED_19), .b(D_5), .O(ED_25) );
and2 gate( .a(ED_20), .b(D_5_NOT), .O(ED_23) );
and2 gate( .a(ED_21), .b(D_5), .O(ED_22) );
or2  gate( .a(ED_22), .b(ED_23), .O(ED_24) );
or2  gate( .a(ED_24), .b(ED_25), .O(ED_26) );
or2  gate( .a(ED_27), .b(ED_26), .O(N372_OBF);
inv1 gate( .a(D_6), .O(D_6_NOT) );
inv1 gate( .a(D_7), .O(D_7_NOT) );
inv1 gate( .a(N17), .O(N17_NOT) );
and2 gate( .a(N17), .b(D_6_NOT), .O(ED_27) );
and2 gate( .a(N17_NOT), .b(D_6_NOT), .O(ED_28) );
and2 gate( .a(CONST1), .b(D_6), .O(ED_29) );
and2 gate( .a(CONST0), .b(D_6), .O(ED_30) );
and2 gate( .a(ED_27), .b(D_7_NOT), .O(ED_36) );
and2 gate( .a(ED_28), .b(D_7), .O(ED_34) );
and2 gate( .a(ED_29), .b(D_7_NOT), .O(ED_32) );
and2 gate( .a(ED_30), .b(D_7), .O(ED_31) );
or2  gate( .a(ED_31), .b(ED_32), .O(ED_33) );
or2  gate( .a(ED_33), .b(ED_34), .O(ED_35) );
or2  gate( .a(ED_36), .b(ED_35), .O(N17_OBF);
inv1 gate( .a(D_8), .O(D_8_NOT) );
inv1 gate( .a(D_9), .O(D_9_NOT) );
inv1 gate( .a(N381), .O(N381_NOT) );
and2 gate( .a(N381), .b(D_8_NOT), .O(ED_36) );
and2 gate( .a(N381_NOT), .b(D_8_NOT), .O(ED_37) );
and2 gate( .a(CONST1), .b(D_8), .O(ED_38) );
and2 gate( .a(CONST0), .b(D_8), .O(ED_39) );
and2 gate( .a(ED_36), .b(D_9_NOT), .O(ED_45) );
and2 gate( .a(ED_37), .b(D_9), .O(ED_43) );
and2 gate( .a(ED_38), .b(D_9_NOT), .O(ED_41) );
and2 gate( .a(ED_39), .b(D_9), .O(ED_40) );
or2  gate( .a(ED_40), .b(ED_41), .O(ED_42) );
or2  gate( .a(ED_42), .b(ED_43), .O(ED_44) );
or2  gate( .a(ED_45), .b(ED_44), .O(N381_OBF);
inv1 gate( .a(D_10), .O(D_10_NOT) );
inv1 gate( .a(D_11), .O(D_11_NOT) );
inv1 gate( .a(N381), .O(N381_NOT) );
and2 gate( .a(N381), .b(D_10_NOT), .O(ED_45) );
and2 gate( .a(N381_NOT), .b(D_10_NOT), .O(ED_46) );
and2 gate( .a(CONST1), .b(D_10), .O(ED_47) );
and2 gate( .a(CONST0), .b(D_10), .O(ED_48) );
and2 gate( .a(ED_45), .b(D_11_NOT), .O(ED_54) );
and2 gate( .a(ED_46), .b(D_11), .O(ED_52) );
and2 gate( .a(ED_47), .b(D_11_NOT), .O(ED_50) );
and2 gate( .a(ED_48), .b(D_11), .O(ED_49) );
or2  gate( .a(ED_49), .b(ED_50), .O(ED_51) );
or2  gate( .a(ED_51), .b(ED_52), .O(ED_53) );
or2  gate( .a(ED_54), .b(ED_53), .O(N381_OBF);
inv1 gate( .a(D_12), .O(D_12_NOT) );
inv1 gate( .a(D_13), .O(D_13_NOT) );
inv1 gate( .a(N386), .O(N386_NOT) );
and2 gate( .a(N386), .b(D_12_NOT), .O(ED_54) );
and2 gate( .a(N386_NOT), .b(D_12_NOT), .O(ED_55) );
and2 gate( .a(CONST1), .b(D_12), .O(ED_56) );
and2 gate( .a(CONST0), .b(D_12), .O(ED_57) );
and2 gate( .a(ED_54), .b(D_13_NOT), .O(ED_63) );
and2 gate( .a(ED_55), .b(D_13), .O(ED_61) );
and2 gate( .a(ED_56), .b(D_13_NOT), .O(ED_59) );
and2 gate( .a(ED_57), .b(D_13), .O(ED_58) );
or2  gate( .a(ED_58), .b(ED_59), .O(ED_60) );
or2  gate( .a(ED_60), .b(ED_61), .O(ED_62) );
or2  gate( .a(ED_63), .b(ED_62), .O(N386_OBF);
inv1 gate( .a(D_14), .O(D_14_NOT) );
inv1 gate( .a(D_15), .O(D_15_NOT) );
inv1 gate( .a(N422), .O(N422_NOT) );
and2 gate( .a(N422), .b(D_14_NOT), .O(ED_63) );
and2 gate( .a(N422_NOT), .b(D_14_NOT), .O(ED_64) );
and2 gate( .a(CONST1), .b(D_14), .O(ED_65) );
and2 gate( .a(CONST0), .b(D_14), .O(ED_66) );
and2 gate( .a(ED_63), .b(D_15_NOT), .O(ED_72) );
and2 gate( .a(ED_64), .b(D_15), .O(ED_70) );
and2 gate( .a(ED_65), .b(D_15_NOT), .O(ED_68) );
and2 gate( .a(ED_66), .b(D_15), .O(ED_67) );
or2  gate( .a(ED_67), .b(ED_68), .O(ED_69) );
or2  gate( .a(ED_69), .b(ED_70), .O(ED_71) );
or2  gate( .a(ED_72), .b(ED_71), .O(N422_OBF);
inv1 gate( .a(D_16), .O(D_16_NOT) );
inv1 gate( .a(D_17), .O(D_17_NOT) );
inv1 gate( .a(N399), .O(N399_NOT) );
and2 gate( .a(N399), .b(D_16_NOT), .O(ED_72) );
and2 gate( .a(N399_NOT), .b(D_16_NOT), .O(ED_73) );
and2 gate( .a(CONST1), .b(D_16), .O(ED_74) );
and2 gate( .a(CONST0), .b(D_16), .O(ED_75) );
and2 gate( .a(ED_72), .b(D_17_NOT), .O(ED_81) );
and2 gate( .a(ED_73), .b(D_17), .O(ED_79) );
and2 gate( .a(ED_74), .b(D_17_NOT), .O(ED_77) );
and2 gate( .a(ED_75), .b(D_17), .O(ED_76) );
or2  gate( .a(ED_76), .b(ED_77), .O(ED_78) );
or2  gate( .a(ED_78), .b(ED_79), .O(ED_80) );
or2  gate( .a(ED_81), .b(ED_80), .O(N399_OBF);
inv1 gate( .a(D_18), .O(D_18_NOT) );
inv1 gate( .a(D_19), .O(D_19_NOT) );
inv1 gate( .a(N430), .O(N430_NOT) );
and2 gate( .a(N430), .b(D_18_NOT), .O(ED_81) );
and2 gate( .a(N430_NOT), .b(D_18_NOT), .O(ED_82) );
and2 gate( .a(CONST1), .b(D_18), .O(ED_83) );
and2 gate( .a(CONST0), .b(D_18), .O(ED_84) );
and2 gate( .a(ED_81), .b(D_19_NOT), .O(ED_90) );
and2 gate( .a(ED_82), .b(D_19), .O(ED_88) );
and2 gate( .a(ED_83), .b(D_19_NOT), .O(ED_86) );
and2 gate( .a(ED_84), .b(D_19), .O(ED_85) );
or2  gate( .a(ED_85), .b(ED_86), .O(ED_87) );
or2  gate( .a(ED_87), .b(ED_88), .O(ED_89) );
or2  gate( .a(ED_90), .b(ED_89), .O(N430_OBF);

endmodule
