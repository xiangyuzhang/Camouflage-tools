
module c432 (N1, NO);

input N1;

output NO;

wire ;

inv1 gate1( .a(N1), .O(NO) );


endmodule