
module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);

input  N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,      N99,N102,N105,N108,N112,N115,CONST1,CONST0 //RE__PI;

input D_0,D_1,D_2,D_3,D_4,D_5,D_6,D_7,D_8,D_9,D_10,D_11,D_12,D_13,D_14,D_15,D_16,D_17,D_18,D_19,D_20,D_21,D_22,D_23,D_24,D_25,D_26,D_27,D_28,D_29,D_30,D_31,D_32,D_33,D_34,D_35,D_36,D_37,D_38,D_39,D_40,D_41,D_42,D_43,D_44,D_45,D_46,D_47,D_48,D_49,D_50,D_51,D_52,D_53,D_54,D_55,D_56,D_57,D_58,D_59,D_60,D_61,D_62,D_63,D_64,D_65,D_66,D_67,D_68,D_69,D_70,D_71,D_72,D_73,D_74,D_75,D_76,D_77,D_78,D_79,D_80,D_81,D_82,D_83,D_84,D_85,D_86,D_87,D_88,D_89,D_90,D_91,D_92,D_93,D_94,D_95,D_96,D_97,D_98,D_99 //RE__ALLOW(00,01,10,11);

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429,D_0_NOT,D_1_NOT,N246_NOT,N246_OBF,ED_0,ED_1,ED_2,ED_3,ED_4,ED_5,ED_6,ED_7,ED_8,ED_9,D_2_NOT,D_3_NOT,N336_NOT,N336_OBF,ED_9,ED_10,ED_11,ED_12,ED_13,ED_14,ED_15,ED_16,ED_17,ED_18,D_4_NOT,D_5_NOT,N372_NOT,N372_OBF,ED_18,ED_19,ED_20,ED_21,ED_22,ED_23,ED_24,ED_25,ED_26,ED_27,D_6_NOT,D_7_NOT,N17_NOT,N17_OBF,ED_27,ED_28,ED_29,ED_30,ED_31,ED_32,ED_33,ED_34,ED_35,ED_36,D_8_NOT,D_9_NOT,N381_NOT,N381_OBF,ED_36,ED_37,ED_38,ED_39,ED_40,ED_41,ED_42,ED_43,ED_44,ED_45,D_10_NOT,D_11_NOT,N381_NOT,N381_OBF,ED_45,ED_46,ED_47,ED_48,ED_49,ED_50,ED_51,ED_52,ED_53,ED_54,D_12_NOT,D_13_NOT,N386_NOT,N386_OBF,ED_54,ED_55,ED_56,ED_57,ED_58,ED_59,ED_60,ED_61,ED_62,ED_63,D_14_NOT,D_15_NOT,N422_NOT,N422_OBF,ED_63,ED_64,ED_65,ED_66,ED_67,ED_68,ED_69,ED_70,ED_71,ED_72,D_16_NOT,D_17_NOT,N399_NOT,N399_OBF,ED_72,ED_73,ED_74,ED_75,ED_76,ED_77,ED_78,ED_79,ED_80,ED_81,D_18_NOT,D_19_NOT,N430_NOT,N430_OBF,ED_81,ED_82,ED_83,ED_84,ED_85,ED_86,ED_87,ED_88,ED_89,ED_90,D_20_NOT,D_21_NOT,N386_NOT,N386_OBF,ED_90,ED_91,ED_92,ED_93,ED_94,ED_95,ED_96,ED_97,ED_98,ED_99,D_22_NOT,D_23_NOT,N393_NOT,N393_OBF,ED_99,ED_100,ED_101,ED_102,ED_103,ED_104,ED_105,ED_106,ED_107,ED_108,D_24_NOT,D_25_NOT,N407_NOT,N407_OBF,ED_108,ED_109,ED_110,ED_111,ED_112,ED_113,ED_114,ED_115,ED_116,ED_117,D_26_NOT,D_27_NOT,N420_NOT,N420_OBF,ED_117,ED_118,ED_119,ED_120,ED_121,ED_122,ED_123,ED_124,ED_125,ED_126,D_28_NOT,D_29_NOT,N429_NOT,N429_OBF,ED_126,ED_127,ED_128,ED_129,ED_130,ED_131,ED_132,ED_133,ED_134,ED_135,D_30_NOT,D_31_NOT,N254_NOT,N254_OBF,ED_135,ED_136,ED_137,ED_138,ED_139,ED_140,ED_141,ED_142,ED_143,ED_144,D_32_NOT,D_33_NOT,N340_NOT,N340_OBF,ED_144,ED_145,ED_146,ED_147,ED_148,ED_149,ED_150,ED_151,ED_152,ED_153,D_34_NOT,D_35_NOT,N374_NOT,N374_OBF,ED_153,ED_154,ED_155,ED_156,ED_157,ED_158,ED_159,ED_160,ED_161,ED_162,D_36_NOT,D_37_NOT,N43_NOT,N43_OBF,ED_162,ED_163,ED_164,ED_165,ED_166,ED_167,ED_168,ED_169,ED_170,ED_171,D_38_NOT,D_39_NOT,N393_NOT,N393_OBF,ED_171,ED_172,ED_173,ED_174,ED_175,ED_176,ED_177,ED_178,ED_179,ED_180,D_40_NOT,D_41_NOT,N257_NOT,N257_OBF,ED_180,ED_181,ED_182,ED_183,ED_184,ED_185,ED_186,ED_187,ED_188,ED_189,D_42_NOT,D_43_NOT,N345_NOT,N345_OBF,ED_189,ED_190,ED_191,ED_192,ED_193,ED_194,ED_195,ED_196,ED_197,ED_198,D_44_NOT,D_45_NOT,N377_NOT,N377_OBF,ED_198,ED_199,ED_200,ED_201,ED_202,ED_203,ED_204,ED_205,ED_206,ED_207,D_46_NOT,D_47_NOT,N82_NOT,N82_OBF,ED_207,ED_208,ED_209,ED_210,ED_211,ED_212,ED_213,ED_214,ED_215,ED_216,D_48_NOT,D_49_NOT,N407_NOT,N407_OBF,ED_216,ED_217,ED_218,ED_219,ED_220,ED_221,ED_222,ED_223,ED_224,ED_225,D_50_NOT,D_51_NOT,N386_NOT,N386_OBF,ED_225,ED_226,ED_227,ED_228,ED_229,ED_230,ED_231,ED_232,ED_233,ED_234,D_52_NOT,D_53_NOT,N393_NOT,N393_OBF,ED_234,ED_235,ED_236,ED_237,ED_238,ED_239,ED_240,ED_241,ED_242,ED_243,D_54_NOT,D_55_NOT,N418_NOT,N418_OBF,ED_243,ED_244,ED_245,ED_246,ED_247,ED_248,ED_249,ED_250,ED_251,ED_252,D_56_NOT,D_57_NOT,N399_NOT,N399_OBF,ED_252,ED_253,ED_254,ED_255,ED_256,ED_257,ED_258,ED_259,ED_260,ED_261,D_58_NOT,D_59_NOT,N425_NOT,N425_OBF,ED_261,ED_262,ED_263,ED_264,ED_265,ED_266,ED_267,ED_268,ED_269,ED_270,D_60_NOT,D_61_NOT,N4_NOT,N4_OBF,ED_270,ED_271,ED_272,ED_273,ED_274,ED_275,ED_276,ED_277,ED_278,ED_279,D_62_NOT,D_63_NOT,N242_NOT,N242_OBF,ED_279,ED_280,ED_281,ED_282,ED_283,ED_284,ED_285,ED_286,ED_287,ED_288,D_64_NOT,D_65_NOT,N334_NOT,N334_OBF,ED_288,ED_289,ED_290,ED_291,ED_292,ED_293,ED_294,ED_295,ED_296,ED_297,D_66_NOT,D_67_NOT,N371_NOT,N371_OBF,ED_297,ED_298,ED_299,ED_300,ED_301,ED_302,ED_303,ED_304,ED_305,ED_306,D_68_NOT,D_69_NOT,N380_NOT,N380_OBF,ED_306,ED_307,ED_308,ED_309,ED_310,ED_311,ED_312,ED_313,ED_314,ED_315,D_70_NOT,D_71_NOT,N381_NOT,N381_OBF,ED_315,ED_316,ED_317,ED_318,ED_319,ED_320,ED_321,ED_322,ED_323,ED_324,D_72_NOT,D_73_NOT,N422_NOT,N422_OBF,ED_324,ED_325,ED_326,ED_327,ED_328,ED_329,ED_330,ED_331,ED_332,ED_333,D_74_NOT,D_75_NOT,N425_NOT,N425_OBF,ED_333,ED_334,ED_335,ED_336,ED_337,ED_338,ED_339,ED_340,ED_341,ED_342,D_76_NOT,D_77_NOT,N429_NOT,N429_OBF,ED_342,ED_343,ED_344,ED_345,ED_346,ED_347,ED_348,ED_349,ED_350,ED_351,D_78_NOT,D_79_NOT,N432_NOT,N432_OBF,ED_351,ED_352,ED_353,ED_354,ED_355,ED_356,ED_357,ED_358,ED_359,ED_360,D_80_NOT,D_81_NOT,N381_NOT,N381_OBF,ED_360,ED_361,ED_362,ED_363,ED_364,ED_365,ED_366,ED_367,ED_368,ED_369,D_82_NOT,D_83_NOT,N386_NOT,N386_OBF,ED_369,ED_370,ED_371,ED_372,ED_373,ED_374,ED_375,ED_376,ED_377,ED_378,D_84_NOT,D_85_NOT,N425_NOT,N425_OBF,ED_378,ED_379,ED_380,ED_381,ED_382,ED_383,ED_384,ED_385,ED_386,ED_387,D_86_NOT,D_87_NOT,N428_NOT,N428_OBF,ED_387,ED_388,ED_389,ED_390,ED_391,ED_392,ED_393,ED_394,ED_395,ED_396,D_88_NOT,D_89_NOT,N431_NOT,N431_OBF,ED_396,ED_397,ED_398,ED_399,ED_400,ED_401,ED_402,ED_403,ED_404,ED_405,D_90_NOT,D_91_NOT,N258_NOT,N258_OBF,ED_405,ED_406,ED_407,ED_408,ED_409,ED_410,ED_411,ED_412,ED_413,ED_414,D_92_NOT,D_93_NOT,N346_NOT,N346_OBF,ED_414,ED_415,ED_416,ED_417,ED_418,ED_419,ED_420,ED_421,ED_422,ED_423,D_94_NOT,D_95_NOT,N378_NOT,N378_OBF,ED_423,ED_424,ED_425,ED_426,ED_427,ED_428,ED_429,ED_430,ED_431,ED_432,D_96_NOT,D_97_NOT,N95_NOT,N95_OBF,ED_432,ED_433,ED_434,ED_435,ED_436,ED_437,ED_438,ED_439,ED_440,ED_441,D_98_NOT,D_99_NOT,N411_NOT,N411_OBF,ED_441,ED_442,ED_443,ED_444,ED_445,ED_446,ED_447,ED_448,ED_449,ED_450;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );
nand2 gate78( .a(N227), .b(N184), .O(N288) );
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );
nand2 gate135( .a(N360), .b(N92), .O(N377) );
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4_OBF), .b(N242_OBF), .c(N334_OBF), .d(N371_OBF), .O(N380_OBF) );
nand4 gate139( .a(N246_OBF), .b(N336_OBF), .c(N372_OBF), .d(N17_OBF), .O(N381_OBF) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254_OBF), .b(N340_OBF), .c(N374_OBF), .d(N43_OBF), .O(N393_OBF) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257_OBF), .b(N345_OBF), .c(N377_OBF), .d(N82_OBF), .O(N407_OBF) );
nand4 gate145( .a(N258_OBF), .b(N346_OBF), .c(N378_OBF), .d(N95_OBF), .O(N411_OBF) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380_OBF), .O(N415) );
and8 gate148( .a(N381_OBF), .b(N386), .c(N393_OBF), .d(N399), .e(N404), .f(N407_OBF), .g(N411_OBF), .h(N414), .O(N416) );
inv1 gate149( .a(N393_OBF), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407_OBF), .O(N419) );
inv1 gate152( .a(N411_OBF), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393_OBF), .c(N418), .d(N399), .O(N425_OBF) );
nand3 gate156( .a(N399), .b(N393_OBF), .c(N419), .O(N428) );
nand4 gate157( .a(N386_OBF), .b(N393_OBF), .c(N407_OBF), .d(N420_OBF), .O(N429_OBF) );
nand4 gate158( .a(N381_OBF), .b(N386), .c(N422), .d(N399), .O(N430_OBF) );
nand4 gate159( .a(N381_OBF), .b(N386), .c(N425_OBF), .d(N428), .O(N431_OBF) );
nand4 gate160( .a(N381_OBF), .b(N422), .c(N425_OBF), .d(N429_OBF), .O(N432_OBF) );
inv1 gate( .a(D_0), .O(D_0_NOT) );
inv1 gate( .a(D_1), .O(D_1_NOT) );
inv1 gate( .a(N246), .O(N246_NOT) );
and2 gate( .a(N246), .b(D_0_NOT), .O(ED_0) );
and2 gate( .a(N246_NOT), .b(D_0_NOT), .O(ED_1) );
and2 gate( .a(CONST1), .b(D_0), .O(ED_2) );
and2 gate( .a(CONST0), .b(D_0), .O(ED_3) );
and2 gate( .a(ED_0), .b(D_1_NOT), .O(ED_9) );
and2 gate( .a(ED_1), .b(D_1), .O(ED_7) );
and2 gate( .a(ED_2), .b(D_1_NOT), .O(ED_5) );
and2 gate( .a(ED_3), .b(D_1), .O(ED_4) );
or2  gate( .a(ED_4), .b(ED_5), .O(ED_6) );
or2  gate( .a(ED_6), .b(ED_7), .O(ED_8) );
or2  gate( .a(ED_9), .b(ED_8), .O(N246_OBF);
inv1 gate( .a(D_2), .O(D_2_NOT) );
inv1 gate( .a(D_3), .O(D_3_NOT) );
inv1 gate( .a(N336), .O(N336_NOT) );
and2 gate( .a(N336), .b(D_2_NOT), .O(ED_9) );
and2 gate( .a(N336_NOT), .b(D_2_NOT), .O(ED_10) );
and2 gate( .a(CONST1), .b(D_2), .O(ED_11) );
and2 gate( .a(CONST0), .b(D_2), .O(ED_12) );
and2 gate( .a(ED_9), .b(D_3_NOT), .O(ED_18) );
and2 gate( .a(ED_10), .b(D_3), .O(ED_16) );
and2 gate( .a(ED_11), .b(D_3_NOT), .O(ED_14) );
and2 gate( .a(ED_12), .b(D_3), .O(ED_13) );
or2  gate( .a(ED_13), .b(ED_14), .O(ED_15) );
or2  gate( .a(ED_15), .b(ED_16), .O(ED_17) );
or2  gate( .a(ED_18), .b(ED_17), .O(N336_OBF);
inv1 gate( .a(D_4), .O(D_4_NOT) );
inv1 gate( .a(D_5), .O(D_5_NOT) );
inv1 gate( .a(N372), .O(N372_NOT) );
and2 gate( .a(N372), .b(D_4_NOT), .O(ED_18) );
and2 gate( .a(N372_NOT), .b(D_4_NOT), .O(ED_19) );
and2 gate( .a(CONST1), .b(D_4), .O(ED_20) );
and2 gate( .a(CONST0), .b(D_4), .O(ED_21) );
and2 gate( .a(ED_18), .b(D_5_NOT), .O(ED_27) );
and2 gate( .a(ED_19), .b(D_5), .O(ED_25) );
and2 gate( .a(ED_20), .b(D_5_NOT), .O(ED_23) );
and2 gate( .a(ED_21), .b(D_5), .O(ED_22) );
or2  gate( .a(ED_22), .b(ED_23), .O(ED_24) );
or2  gate( .a(ED_24), .b(ED_25), .O(ED_26) );
or2  gate( .a(ED_27), .b(ED_26), .O(N372_OBF);
inv1 gate( .a(D_6), .O(D_6_NOT) );
inv1 gate( .a(D_7), .O(D_7_NOT) );
inv1 gate( .a(N17), .O(N17_NOT) );
and2 gate( .a(N17), .b(D_6_NOT), .O(ED_27) );
and2 gate( .a(N17_NOT), .b(D_6_NOT), .O(ED_28) );
and2 gate( .a(CONST1), .b(D_6), .O(ED_29) );
and2 gate( .a(CONST0), .b(D_6), .O(ED_30) );
and2 gate( .a(ED_27), .b(D_7_NOT), .O(ED_36) );
and2 gate( .a(ED_28), .b(D_7), .O(ED_34) );
and2 gate( .a(ED_29), .b(D_7_NOT), .O(ED_32) );
and2 gate( .a(ED_30), .b(D_7), .O(ED_31) );
or2  gate( .a(ED_31), .b(ED_32), .O(ED_33) );
or2  gate( .a(ED_33), .b(ED_34), .O(ED_35) );
or2  gate( .a(ED_36), .b(ED_35), .O(N17_OBF);
inv1 gate( .a(D_8), .O(D_8_NOT) );
inv1 gate( .a(D_9), .O(D_9_NOT) );
inv1 gate( .a(N381), .O(N381_NOT) );
and2 gate( .a(N381), .b(D_8_NOT), .O(ED_36) );
and2 gate( .a(N381_NOT), .b(D_8_NOT), .O(ED_37) );
and2 gate( .a(CONST1), .b(D_8), .O(ED_38) );
and2 gate( .a(CONST0), .b(D_8), .O(ED_39) );
and2 gate( .a(ED_36), .b(D_9_NOT), .O(ED_45) );
and2 gate( .a(ED_37), .b(D_9), .O(ED_43) );
and2 gate( .a(ED_38), .b(D_9_NOT), .O(ED_41) );
and2 gate( .a(ED_39), .b(D_9), .O(ED_40) );
or2  gate( .a(ED_40), .b(ED_41), .O(ED_42) );
or2  gate( .a(ED_42), .b(ED_43), .O(ED_44) );
or2  gate( .a(ED_45), .b(ED_44), .O(N381_OBF);
inv1 gate( .a(D_10), .O(D_10_NOT) );
inv1 gate( .a(D_11), .O(D_11_NOT) );
inv1 gate( .a(N381), .O(N381_NOT) );
and2 gate( .a(N381), .b(D_10_NOT), .O(ED_45) );
and2 gate( .a(N381_NOT), .b(D_10_NOT), .O(ED_46) );
and2 gate( .a(CONST1), .b(D_10), .O(ED_47) );
and2 gate( .a(CONST0), .b(D_10), .O(ED_48) );
and2 gate( .a(ED_45), .b(D_11_NOT), .O(ED_54) );
and2 gate( .a(ED_46), .b(D_11), .O(ED_52) );
and2 gate( .a(ED_47), .b(D_11_NOT), .O(ED_50) );
and2 gate( .a(ED_48), .b(D_11), .O(ED_49) );
or2  gate( .a(ED_49), .b(ED_50), .O(ED_51) );
or2  gate( .a(ED_51), .b(ED_52), .O(ED_53) );
or2  gate( .a(ED_54), .b(ED_53), .O(N381_OBF);
inv1 gate( .a(D_12), .O(D_12_NOT) );
inv1 gate( .a(D_13), .O(D_13_NOT) );
inv1 gate( .a(N386), .O(N386_NOT) );
and2 gate( .a(N386), .b(D_12_NOT), .O(ED_54) );
and2 gate( .a(N386_NOT), .b(D_12_NOT), .O(ED_55) );
and2 gate( .a(CONST1), .b(D_12), .O(ED_56) );
and2 gate( .a(CONST0), .b(D_12), .O(ED_57) );
and2 gate( .a(ED_54), .b(D_13_NOT), .O(ED_63) );
and2 gate( .a(ED_55), .b(D_13), .O(ED_61) );
and2 gate( .a(ED_56), .b(D_13_NOT), .O(ED_59) );
and2 gate( .a(ED_57), .b(D_13), .O(ED_58) );
or2  gate( .a(ED_58), .b(ED_59), .O(ED_60) );
or2  gate( .a(ED_60), .b(ED_61), .O(ED_62) );
or2  gate( .a(ED_63), .b(ED_62), .O(N386_OBF);
inv1 gate( .a(D_14), .O(D_14_NOT) );
inv1 gate( .a(D_15), .O(D_15_NOT) );
inv1 gate( .a(N422), .O(N422_NOT) );
and2 gate( .a(N422), .b(D_14_NOT), .O(ED_63) );
and2 gate( .a(N422_NOT), .b(D_14_NOT), .O(ED_64) );
and2 gate( .a(CONST1), .b(D_14), .O(ED_65) );
and2 gate( .a(CONST0), .b(D_14), .O(ED_66) );
and2 gate( .a(ED_63), .b(D_15_NOT), .O(ED_72) );
and2 gate( .a(ED_64), .b(D_15), .O(ED_70) );
and2 gate( .a(ED_65), .b(D_15_NOT), .O(ED_68) );
and2 gate( .a(ED_66), .b(D_15), .O(ED_67) );
or2  gate( .a(ED_67), .b(ED_68), .O(ED_69) );
or2  gate( .a(ED_69), .b(ED_70), .O(ED_71) );
or2  gate( .a(ED_72), .b(ED_71), .O(N422_OBF);
inv1 gate( .a(D_16), .O(D_16_NOT) );
inv1 gate( .a(D_17), .O(D_17_NOT) );
inv1 gate( .a(N399), .O(N399_NOT) );
and2 gate( .a(N399), .b(D_16_NOT), .O(ED_72) );
and2 gate( .a(N399_NOT), .b(D_16_NOT), .O(ED_73) );
and2 gate( .a(CONST1), .b(D_16), .O(ED_74) );
and2 gate( .a(CONST0), .b(D_16), .O(ED_75) );
and2 gate( .a(ED_72), .b(D_17_NOT), .O(ED_81) );
and2 gate( .a(ED_73), .b(D_17), .O(ED_79) );
and2 gate( .a(ED_74), .b(D_17_NOT), .O(ED_77) );
and2 gate( .a(ED_75), .b(D_17), .O(ED_76) );
or2  gate( .a(ED_76), .b(ED_77), .O(ED_78) );
or2  gate( .a(ED_78), .b(ED_79), .O(ED_80) );
or2  gate( .a(ED_81), .b(ED_80), .O(N399_OBF);
inv1 gate( .a(D_18), .O(D_18_NOT) );
inv1 gate( .a(D_19), .O(D_19_NOT) );
inv1 gate( .a(N430), .O(N430_NOT) );
and2 gate( .a(N430), .b(D_18_NOT), .O(ED_81) );
and2 gate( .a(N430_NOT), .b(D_18_NOT), .O(ED_82) );
and2 gate( .a(CONST1), .b(D_18), .O(ED_83) );
and2 gate( .a(CONST0), .b(D_18), .O(ED_84) );
and2 gate( .a(ED_81), .b(D_19_NOT), .O(ED_90) );
and2 gate( .a(ED_82), .b(D_19), .O(ED_88) );
and2 gate( .a(ED_83), .b(D_19_NOT), .O(ED_86) );
and2 gate( .a(ED_84), .b(D_19), .O(ED_85) );
or2  gate( .a(ED_85), .b(ED_86), .O(ED_87) );
or2  gate( .a(ED_87), .b(ED_88), .O(ED_89) );
or2  gate( .a(ED_90), .b(ED_89), .O(N430_OBF);
inv1 gate( .a(D_20), .O(D_20_NOT) );
inv1 gate( .a(D_21), .O(D_21_NOT) );
inv1 gate( .a(N386), .O(N386_NOT) );
and2 gate( .a(N386), .b(D_20_NOT), .O(ED_90) );
and2 gate( .a(N386_NOT), .b(D_20_NOT), .O(ED_91) );
and2 gate( .a(CONST1), .b(D_20), .O(ED_92) );
and2 gate( .a(CONST0), .b(D_20), .O(ED_93) );
and2 gate( .a(ED_90), .b(D_21_NOT), .O(ED_99) );
and2 gate( .a(ED_91), .b(D_21), .O(ED_97) );
and2 gate( .a(ED_92), .b(D_21_NOT), .O(ED_95) );
and2 gate( .a(ED_93), .b(D_21), .O(ED_94) );
or2  gate( .a(ED_94), .b(ED_95), .O(ED_96) );
or2  gate( .a(ED_96), .b(ED_97), .O(ED_98) );
or2  gate( .a(ED_99), .b(ED_98), .O(N386_OBF);
inv1 gate( .a(D_22), .O(D_22_NOT) );
inv1 gate( .a(D_23), .O(D_23_NOT) );
inv1 gate( .a(N393), .O(N393_NOT) );
and2 gate( .a(N393), .b(D_22_NOT), .O(ED_99) );
and2 gate( .a(N393_NOT), .b(D_22_NOT), .O(ED_100) );
and2 gate( .a(CONST1), .b(D_22), .O(ED_101) );
and2 gate( .a(CONST0), .b(D_22), .O(ED_102) );
and2 gate( .a(ED_99), .b(D_23_NOT), .O(ED_108) );
and2 gate( .a(ED_100), .b(D_23), .O(ED_106) );
and2 gate( .a(ED_101), .b(D_23_NOT), .O(ED_104) );
and2 gate( .a(ED_102), .b(D_23), .O(ED_103) );
or2  gate( .a(ED_103), .b(ED_104), .O(ED_105) );
or2  gate( .a(ED_105), .b(ED_106), .O(ED_107) );
or2  gate( .a(ED_108), .b(ED_107), .O(N393_OBF);
inv1 gate( .a(D_24), .O(D_24_NOT) );
inv1 gate( .a(D_25), .O(D_25_NOT) );
inv1 gate( .a(N407), .O(N407_NOT) );
and2 gate( .a(N407), .b(D_24_NOT), .O(ED_108) );
and2 gate( .a(N407_NOT), .b(D_24_NOT), .O(ED_109) );
and2 gate( .a(CONST1), .b(D_24), .O(ED_110) );
and2 gate( .a(CONST0), .b(D_24), .O(ED_111) );
and2 gate( .a(ED_108), .b(D_25_NOT), .O(ED_117) );
and2 gate( .a(ED_109), .b(D_25), .O(ED_115) );
and2 gate( .a(ED_110), .b(D_25_NOT), .O(ED_113) );
and2 gate( .a(ED_111), .b(D_25), .O(ED_112) );
or2  gate( .a(ED_112), .b(ED_113), .O(ED_114) );
or2  gate( .a(ED_114), .b(ED_115), .O(ED_116) );
or2  gate( .a(ED_117), .b(ED_116), .O(N407_OBF);
inv1 gate( .a(D_26), .O(D_26_NOT) );
inv1 gate( .a(D_27), .O(D_27_NOT) );
inv1 gate( .a(N420), .O(N420_NOT) );
and2 gate( .a(N420), .b(D_26_NOT), .O(ED_117) );
and2 gate( .a(N420_NOT), .b(D_26_NOT), .O(ED_118) );
and2 gate( .a(CONST1), .b(D_26), .O(ED_119) );
and2 gate( .a(CONST0), .b(D_26), .O(ED_120) );
and2 gate( .a(ED_117), .b(D_27_NOT), .O(ED_126) );
and2 gate( .a(ED_118), .b(D_27), .O(ED_124) );
and2 gate( .a(ED_119), .b(D_27_NOT), .O(ED_122) );
and2 gate( .a(ED_120), .b(D_27), .O(ED_121) );
or2  gate( .a(ED_121), .b(ED_122), .O(ED_123) );
or2  gate( .a(ED_123), .b(ED_124), .O(ED_125) );
or2  gate( .a(ED_126), .b(ED_125), .O(N420_OBF);
inv1 gate( .a(D_28), .O(D_28_NOT) );
inv1 gate( .a(D_29), .O(D_29_NOT) );
inv1 gate( .a(N429), .O(N429_NOT) );
and2 gate( .a(N429), .b(D_28_NOT), .O(ED_126) );
and2 gate( .a(N429_NOT), .b(D_28_NOT), .O(ED_127) );
and2 gate( .a(CONST1), .b(D_28), .O(ED_128) );
and2 gate( .a(CONST0), .b(D_28), .O(ED_129) );
and2 gate( .a(ED_126), .b(D_29_NOT), .O(ED_135) );
and2 gate( .a(ED_127), .b(D_29), .O(ED_133) );
and2 gate( .a(ED_128), .b(D_29_NOT), .O(ED_131) );
and2 gate( .a(ED_129), .b(D_29), .O(ED_130) );
or2  gate( .a(ED_130), .b(ED_131), .O(ED_132) );
or2  gate( .a(ED_132), .b(ED_133), .O(ED_134) );
or2  gate( .a(ED_135), .b(ED_134), .O(N429_OBF);
inv1 gate( .a(D_30), .O(D_30_NOT) );
inv1 gate( .a(D_31), .O(D_31_NOT) );
inv1 gate( .a(N254), .O(N254_NOT) );
and2 gate( .a(N254), .b(D_30_NOT), .O(ED_135) );
and2 gate( .a(N254_NOT), .b(D_30_NOT), .O(ED_136) );
and2 gate( .a(CONST1), .b(D_30), .O(ED_137) );
and2 gate( .a(CONST0), .b(D_30), .O(ED_138) );
and2 gate( .a(ED_135), .b(D_31_NOT), .O(ED_144) );
and2 gate( .a(ED_136), .b(D_31), .O(ED_142) );
and2 gate( .a(ED_137), .b(D_31_NOT), .O(ED_140) );
and2 gate( .a(ED_138), .b(D_31), .O(ED_139) );
or2  gate( .a(ED_139), .b(ED_140), .O(ED_141) );
or2  gate( .a(ED_141), .b(ED_142), .O(ED_143) );
or2  gate( .a(ED_144), .b(ED_143), .O(N254_OBF);
inv1 gate( .a(D_32), .O(D_32_NOT) );
inv1 gate( .a(D_33), .O(D_33_NOT) );
inv1 gate( .a(N340), .O(N340_NOT) );
and2 gate( .a(N340), .b(D_32_NOT), .O(ED_144) );
and2 gate( .a(N340_NOT), .b(D_32_NOT), .O(ED_145) );
and2 gate( .a(CONST1), .b(D_32), .O(ED_146) );
and2 gate( .a(CONST0), .b(D_32), .O(ED_147) );
and2 gate( .a(ED_144), .b(D_33_NOT), .O(ED_153) );
and2 gate( .a(ED_145), .b(D_33), .O(ED_151) );
and2 gate( .a(ED_146), .b(D_33_NOT), .O(ED_149) );
and2 gate( .a(ED_147), .b(D_33), .O(ED_148) );
or2  gate( .a(ED_148), .b(ED_149), .O(ED_150) );
or2  gate( .a(ED_150), .b(ED_151), .O(ED_152) );
or2  gate( .a(ED_153), .b(ED_152), .O(N340_OBF);
inv1 gate( .a(D_34), .O(D_34_NOT) );
inv1 gate( .a(D_35), .O(D_35_NOT) );
inv1 gate( .a(N374), .O(N374_NOT) );
and2 gate( .a(N374), .b(D_34_NOT), .O(ED_153) );
and2 gate( .a(N374_NOT), .b(D_34_NOT), .O(ED_154) );
and2 gate( .a(CONST1), .b(D_34), .O(ED_155) );
and2 gate( .a(CONST0), .b(D_34), .O(ED_156) );
and2 gate( .a(ED_153), .b(D_35_NOT), .O(ED_162) );
and2 gate( .a(ED_154), .b(D_35), .O(ED_160) );
and2 gate( .a(ED_155), .b(D_35_NOT), .O(ED_158) );
and2 gate( .a(ED_156), .b(D_35), .O(ED_157) );
or2  gate( .a(ED_157), .b(ED_158), .O(ED_159) );
or2  gate( .a(ED_159), .b(ED_160), .O(ED_161) );
or2  gate( .a(ED_162), .b(ED_161), .O(N374_OBF);
inv1 gate( .a(D_36), .O(D_36_NOT) );
inv1 gate( .a(D_37), .O(D_37_NOT) );
inv1 gate( .a(N43), .O(N43_NOT) );
and2 gate( .a(N43), .b(D_36_NOT), .O(ED_162) );
and2 gate( .a(N43_NOT), .b(D_36_NOT), .O(ED_163) );
and2 gate( .a(CONST1), .b(D_36), .O(ED_164) );
and2 gate( .a(CONST0), .b(D_36), .O(ED_165) );
and2 gate( .a(ED_162), .b(D_37_NOT), .O(ED_171) );
and2 gate( .a(ED_163), .b(D_37), .O(ED_169) );
and2 gate( .a(ED_164), .b(D_37_NOT), .O(ED_167) );
and2 gate( .a(ED_165), .b(D_37), .O(ED_166) );
or2  gate( .a(ED_166), .b(ED_167), .O(ED_168) );
or2  gate( .a(ED_168), .b(ED_169), .O(ED_170) );
or2  gate( .a(ED_171), .b(ED_170), .O(N43_OBF);
inv1 gate( .a(D_38), .O(D_38_NOT) );
inv1 gate( .a(D_39), .O(D_39_NOT) );
inv1 gate( .a(N393), .O(N393_NOT) );
and2 gate( .a(N393), .b(D_38_NOT), .O(ED_171) );
and2 gate( .a(N393_NOT), .b(D_38_NOT), .O(ED_172) );
and2 gate( .a(CONST1), .b(D_38), .O(ED_173) );
and2 gate( .a(CONST0), .b(D_38), .O(ED_174) );
and2 gate( .a(ED_171), .b(D_39_NOT), .O(ED_180) );
and2 gate( .a(ED_172), .b(D_39), .O(ED_178) );
and2 gate( .a(ED_173), .b(D_39_NOT), .O(ED_176) );
and2 gate( .a(ED_174), .b(D_39), .O(ED_175) );
or2  gate( .a(ED_175), .b(ED_176), .O(ED_177) );
or2  gate( .a(ED_177), .b(ED_178), .O(ED_179) );
or2  gate( .a(ED_180), .b(ED_179), .O(N393_OBF);
inv1 gate( .a(D_40), .O(D_40_NOT) );
inv1 gate( .a(D_41), .O(D_41_NOT) );
inv1 gate( .a(N257), .O(N257_NOT) );
and2 gate( .a(N257), .b(D_40_NOT), .O(ED_180) );
and2 gate( .a(N257_NOT), .b(D_40_NOT), .O(ED_181) );
and2 gate( .a(CONST1), .b(D_40), .O(ED_182) );
and2 gate( .a(CONST0), .b(D_40), .O(ED_183) );
and2 gate( .a(ED_180), .b(D_41_NOT), .O(ED_189) );
and2 gate( .a(ED_181), .b(D_41), .O(ED_187) );
and2 gate( .a(ED_182), .b(D_41_NOT), .O(ED_185) );
and2 gate( .a(ED_183), .b(D_41), .O(ED_184) );
or2  gate( .a(ED_184), .b(ED_185), .O(ED_186) );
or2  gate( .a(ED_186), .b(ED_187), .O(ED_188) );
or2  gate( .a(ED_189), .b(ED_188), .O(N257_OBF);
inv1 gate( .a(D_42), .O(D_42_NOT) );
inv1 gate( .a(D_43), .O(D_43_NOT) );
inv1 gate( .a(N345), .O(N345_NOT) );
and2 gate( .a(N345), .b(D_42_NOT), .O(ED_189) );
and2 gate( .a(N345_NOT), .b(D_42_NOT), .O(ED_190) );
and2 gate( .a(CONST1), .b(D_42), .O(ED_191) );
and2 gate( .a(CONST0), .b(D_42), .O(ED_192) );
and2 gate( .a(ED_189), .b(D_43_NOT), .O(ED_198) );
and2 gate( .a(ED_190), .b(D_43), .O(ED_196) );
and2 gate( .a(ED_191), .b(D_43_NOT), .O(ED_194) );
and2 gate( .a(ED_192), .b(D_43), .O(ED_193) );
or2  gate( .a(ED_193), .b(ED_194), .O(ED_195) );
or2  gate( .a(ED_195), .b(ED_196), .O(ED_197) );
or2  gate( .a(ED_198), .b(ED_197), .O(N345_OBF);
inv1 gate( .a(D_44), .O(D_44_NOT) );
inv1 gate( .a(D_45), .O(D_45_NOT) );
inv1 gate( .a(N377), .O(N377_NOT) );
and2 gate( .a(N377), .b(D_44_NOT), .O(ED_198) );
and2 gate( .a(N377_NOT), .b(D_44_NOT), .O(ED_199) );
and2 gate( .a(CONST1), .b(D_44), .O(ED_200) );
and2 gate( .a(CONST0), .b(D_44), .O(ED_201) );
and2 gate( .a(ED_198), .b(D_45_NOT), .O(ED_207) );
and2 gate( .a(ED_199), .b(D_45), .O(ED_205) );
and2 gate( .a(ED_200), .b(D_45_NOT), .O(ED_203) );
and2 gate( .a(ED_201), .b(D_45), .O(ED_202) );
or2  gate( .a(ED_202), .b(ED_203), .O(ED_204) );
or2  gate( .a(ED_204), .b(ED_205), .O(ED_206) );
or2  gate( .a(ED_207), .b(ED_206), .O(N377_OBF);
inv1 gate( .a(D_46), .O(D_46_NOT) );
inv1 gate( .a(D_47), .O(D_47_NOT) );
inv1 gate( .a(N82), .O(N82_NOT) );
and2 gate( .a(N82), .b(D_46_NOT), .O(ED_207) );
and2 gate( .a(N82_NOT), .b(D_46_NOT), .O(ED_208) );
and2 gate( .a(CONST1), .b(D_46), .O(ED_209) );
and2 gate( .a(CONST0), .b(D_46), .O(ED_210) );
and2 gate( .a(ED_207), .b(D_47_NOT), .O(ED_216) );
and2 gate( .a(ED_208), .b(D_47), .O(ED_214) );
and2 gate( .a(ED_209), .b(D_47_NOT), .O(ED_212) );
and2 gate( .a(ED_210), .b(D_47), .O(ED_211) );
or2  gate( .a(ED_211), .b(ED_212), .O(ED_213) );
or2  gate( .a(ED_213), .b(ED_214), .O(ED_215) );
or2  gate( .a(ED_216), .b(ED_215), .O(N82_OBF);
inv1 gate( .a(D_48), .O(D_48_NOT) );
inv1 gate( .a(D_49), .O(D_49_NOT) );
inv1 gate( .a(N407), .O(N407_NOT) );
and2 gate( .a(N407), .b(D_48_NOT), .O(ED_216) );
and2 gate( .a(N407_NOT), .b(D_48_NOT), .O(ED_217) );
and2 gate( .a(CONST1), .b(D_48), .O(ED_218) );
and2 gate( .a(CONST0), .b(D_48), .O(ED_219) );
and2 gate( .a(ED_216), .b(D_49_NOT), .O(ED_225) );
and2 gate( .a(ED_217), .b(D_49), .O(ED_223) );
and2 gate( .a(ED_218), .b(D_49_NOT), .O(ED_221) );
and2 gate( .a(ED_219), .b(D_49), .O(ED_220) );
or2  gate( .a(ED_220), .b(ED_221), .O(ED_222) );
or2  gate( .a(ED_222), .b(ED_223), .O(ED_224) );
or2  gate( .a(ED_225), .b(ED_224), .O(N407_OBF);
inv1 gate( .a(D_50), .O(D_50_NOT) );
inv1 gate( .a(D_51), .O(D_51_NOT) );
inv1 gate( .a(N386), .O(N386_NOT) );
and2 gate( .a(N386), .b(D_50_NOT), .O(ED_225) );
and2 gate( .a(N386_NOT), .b(D_50_NOT), .O(ED_226) );
and2 gate( .a(CONST1), .b(D_50), .O(ED_227) );
and2 gate( .a(CONST0), .b(D_50), .O(ED_228) );
and2 gate( .a(ED_225), .b(D_51_NOT), .O(ED_234) );
and2 gate( .a(ED_226), .b(D_51), .O(ED_232) );
and2 gate( .a(ED_227), .b(D_51_NOT), .O(ED_230) );
and2 gate( .a(ED_228), .b(D_51), .O(ED_229) );
or2  gate( .a(ED_229), .b(ED_230), .O(ED_231) );
or2  gate( .a(ED_231), .b(ED_232), .O(ED_233) );
or2  gate( .a(ED_234), .b(ED_233), .O(N386_OBF);
inv1 gate( .a(D_52), .O(D_52_NOT) );
inv1 gate( .a(D_53), .O(D_53_NOT) );
inv1 gate( .a(N393), .O(N393_NOT) );
and2 gate( .a(N393), .b(D_52_NOT), .O(ED_234) );
and2 gate( .a(N393_NOT), .b(D_52_NOT), .O(ED_235) );
and2 gate( .a(CONST1), .b(D_52), .O(ED_236) );
and2 gate( .a(CONST0), .b(D_52), .O(ED_237) );
and2 gate( .a(ED_234), .b(D_53_NOT), .O(ED_243) );
and2 gate( .a(ED_235), .b(D_53), .O(ED_241) );
and2 gate( .a(ED_236), .b(D_53_NOT), .O(ED_239) );
and2 gate( .a(ED_237), .b(D_53), .O(ED_238) );
or2  gate( .a(ED_238), .b(ED_239), .O(ED_240) );
or2  gate( .a(ED_240), .b(ED_241), .O(ED_242) );
or2  gate( .a(ED_243), .b(ED_242), .O(N393_OBF);
inv1 gate( .a(D_54), .O(D_54_NOT) );
inv1 gate( .a(D_55), .O(D_55_NOT) );
inv1 gate( .a(N418), .O(N418_NOT) );
and2 gate( .a(N418), .b(D_54_NOT), .O(ED_243) );
and2 gate( .a(N418_NOT), .b(D_54_NOT), .O(ED_244) );
and2 gate( .a(CONST1), .b(D_54), .O(ED_245) );
and2 gate( .a(CONST0), .b(D_54), .O(ED_246) );
and2 gate( .a(ED_243), .b(D_55_NOT), .O(ED_252) );
and2 gate( .a(ED_244), .b(D_55), .O(ED_250) );
and2 gate( .a(ED_245), .b(D_55_NOT), .O(ED_248) );
and2 gate( .a(ED_246), .b(D_55), .O(ED_247) );
or2  gate( .a(ED_247), .b(ED_248), .O(ED_249) );
or2  gate( .a(ED_249), .b(ED_250), .O(ED_251) );
or2  gate( .a(ED_252), .b(ED_251), .O(N418_OBF);
inv1 gate( .a(D_56), .O(D_56_NOT) );
inv1 gate( .a(D_57), .O(D_57_NOT) );
inv1 gate( .a(N399), .O(N399_NOT) );
and2 gate( .a(N399), .b(D_56_NOT), .O(ED_252) );
and2 gate( .a(N399_NOT), .b(D_56_NOT), .O(ED_253) );
and2 gate( .a(CONST1), .b(D_56), .O(ED_254) );
and2 gate( .a(CONST0), .b(D_56), .O(ED_255) );
and2 gate( .a(ED_252), .b(D_57_NOT), .O(ED_261) );
and2 gate( .a(ED_253), .b(D_57), .O(ED_259) );
and2 gate( .a(ED_254), .b(D_57_NOT), .O(ED_257) );
and2 gate( .a(ED_255), .b(D_57), .O(ED_256) );
or2  gate( .a(ED_256), .b(ED_257), .O(ED_258) );
or2  gate( .a(ED_258), .b(ED_259), .O(ED_260) );
or2  gate( .a(ED_261), .b(ED_260), .O(N399_OBF);
inv1 gate( .a(D_58), .O(D_58_NOT) );
inv1 gate( .a(D_59), .O(D_59_NOT) );
inv1 gate( .a(N425), .O(N425_NOT) );
and2 gate( .a(N425), .b(D_58_NOT), .O(ED_261) );
and2 gate( .a(N425_NOT), .b(D_58_NOT), .O(ED_262) );
and2 gate( .a(CONST1), .b(D_58), .O(ED_263) );
and2 gate( .a(CONST0), .b(D_58), .O(ED_264) );
and2 gate( .a(ED_261), .b(D_59_NOT), .O(ED_270) );
and2 gate( .a(ED_262), .b(D_59), .O(ED_268) );
and2 gate( .a(ED_263), .b(D_59_NOT), .O(ED_266) );
and2 gate( .a(ED_264), .b(D_59), .O(ED_265) );
or2  gate( .a(ED_265), .b(ED_266), .O(ED_267) );
or2  gate( .a(ED_267), .b(ED_268), .O(ED_269) );
or2  gate( .a(ED_270), .b(ED_269), .O(N425_OBF);
inv1 gate( .a(D_60), .O(D_60_NOT) );
inv1 gate( .a(D_61), .O(D_61_NOT) );
inv1 gate( .a(N4), .O(N4_NOT) );
and2 gate( .a(N4), .b(D_60_NOT), .O(ED_270) );
and2 gate( .a(N4_NOT), .b(D_60_NOT), .O(ED_271) );
and2 gate( .a(CONST1), .b(D_60), .O(ED_272) );
and2 gate( .a(CONST0), .b(D_60), .O(ED_273) );
and2 gate( .a(ED_270), .b(D_61_NOT), .O(ED_279) );
and2 gate( .a(ED_271), .b(D_61), .O(ED_277) );
and2 gate( .a(ED_272), .b(D_61_NOT), .O(ED_275) );
and2 gate( .a(ED_273), .b(D_61), .O(ED_274) );
or2  gate( .a(ED_274), .b(ED_275), .O(ED_276) );
or2  gate( .a(ED_276), .b(ED_277), .O(ED_278) );
or2  gate( .a(ED_279), .b(ED_278), .O(N4_OBF);
inv1 gate( .a(D_62), .O(D_62_NOT) );
inv1 gate( .a(D_63), .O(D_63_NOT) );
inv1 gate( .a(N242), .O(N242_NOT) );
and2 gate( .a(N242), .b(D_62_NOT), .O(ED_279) );
and2 gate( .a(N242_NOT), .b(D_62_NOT), .O(ED_280) );
and2 gate( .a(CONST1), .b(D_62), .O(ED_281) );
and2 gate( .a(CONST0), .b(D_62), .O(ED_282) );
and2 gate( .a(ED_279), .b(D_63_NOT), .O(ED_288) );
and2 gate( .a(ED_280), .b(D_63), .O(ED_286) );
and2 gate( .a(ED_281), .b(D_63_NOT), .O(ED_284) );
and2 gate( .a(ED_282), .b(D_63), .O(ED_283) );
or2  gate( .a(ED_283), .b(ED_284), .O(ED_285) );
or2  gate( .a(ED_285), .b(ED_286), .O(ED_287) );
or2  gate( .a(ED_288), .b(ED_287), .O(N242_OBF);
inv1 gate( .a(D_64), .O(D_64_NOT) );
inv1 gate( .a(D_65), .O(D_65_NOT) );
inv1 gate( .a(N334), .O(N334_NOT) );
and2 gate( .a(N334), .b(D_64_NOT), .O(ED_288) );
and2 gate( .a(N334_NOT), .b(D_64_NOT), .O(ED_289) );
and2 gate( .a(CONST1), .b(D_64), .O(ED_290) );
and2 gate( .a(CONST0), .b(D_64), .O(ED_291) );
and2 gate( .a(ED_288), .b(D_65_NOT), .O(ED_297) );
and2 gate( .a(ED_289), .b(D_65), .O(ED_295) );
and2 gate( .a(ED_290), .b(D_65_NOT), .O(ED_293) );
and2 gate( .a(ED_291), .b(D_65), .O(ED_292) );
or2  gate( .a(ED_292), .b(ED_293), .O(ED_294) );
or2  gate( .a(ED_294), .b(ED_295), .O(ED_296) );
or2  gate( .a(ED_297), .b(ED_296), .O(N334_OBF);
inv1 gate( .a(D_66), .O(D_66_NOT) );
inv1 gate( .a(D_67), .O(D_67_NOT) );
inv1 gate( .a(N371), .O(N371_NOT) );
and2 gate( .a(N371), .b(D_66_NOT), .O(ED_297) );
and2 gate( .a(N371_NOT), .b(D_66_NOT), .O(ED_298) );
and2 gate( .a(CONST1), .b(D_66), .O(ED_299) );
and2 gate( .a(CONST0), .b(D_66), .O(ED_300) );
and2 gate( .a(ED_297), .b(D_67_NOT), .O(ED_306) );
and2 gate( .a(ED_298), .b(D_67), .O(ED_304) );
and2 gate( .a(ED_299), .b(D_67_NOT), .O(ED_302) );
and2 gate( .a(ED_300), .b(D_67), .O(ED_301) );
or2  gate( .a(ED_301), .b(ED_302), .O(ED_303) );
or2  gate( .a(ED_303), .b(ED_304), .O(ED_305) );
or2  gate( .a(ED_306), .b(ED_305), .O(N371_OBF);
inv1 gate( .a(D_68), .O(D_68_NOT) );
inv1 gate( .a(D_69), .O(D_69_NOT) );
inv1 gate( .a(N380), .O(N380_NOT) );
and2 gate( .a(N380), .b(D_68_NOT), .O(ED_306) );
and2 gate( .a(N380_NOT), .b(D_68_NOT), .O(ED_307) );
and2 gate( .a(CONST1), .b(D_68), .O(ED_308) );
and2 gate( .a(CONST0), .b(D_68), .O(ED_309) );
and2 gate( .a(ED_306), .b(D_69_NOT), .O(ED_315) );
and2 gate( .a(ED_307), .b(D_69), .O(ED_313) );
and2 gate( .a(ED_308), .b(D_69_NOT), .O(ED_311) );
and2 gate( .a(ED_309), .b(D_69), .O(ED_310) );
or2  gate( .a(ED_310), .b(ED_311), .O(ED_312) );
or2  gate( .a(ED_312), .b(ED_313), .O(ED_314) );
or2  gate( .a(ED_315), .b(ED_314), .O(N380_OBF);
inv1 gate( .a(D_70), .O(D_70_NOT) );
inv1 gate( .a(D_71), .O(D_71_NOT) );
inv1 gate( .a(N381), .O(N381_NOT) );
and2 gate( .a(N381), .b(D_70_NOT), .O(ED_315) );
and2 gate( .a(N381_NOT), .b(D_70_NOT), .O(ED_316) );
and2 gate( .a(CONST1), .b(D_70), .O(ED_317) );
and2 gate( .a(CONST0), .b(D_70), .O(ED_318) );
and2 gate( .a(ED_315), .b(D_71_NOT), .O(ED_324) );
and2 gate( .a(ED_316), .b(D_71), .O(ED_322) );
and2 gate( .a(ED_317), .b(D_71_NOT), .O(ED_320) );
and2 gate( .a(ED_318), .b(D_71), .O(ED_319) );
or2  gate( .a(ED_319), .b(ED_320), .O(ED_321) );
or2  gate( .a(ED_321), .b(ED_322), .O(ED_323) );
or2  gate( .a(ED_324), .b(ED_323), .O(N381_OBF);
inv1 gate( .a(D_72), .O(D_72_NOT) );
inv1 gate( .a(D_73), .O(D_73_NOT) );
inv1 gate( .a(N422), .O(N422_NOT) );
and2 gate( .a(N422), .b(D_72_NOT), .O(ED_324) );
and2 gate( .a(N422_NOT), .b(D_72_NOT), .O(ED_325) );
and2 gate( .a(CONST1), .b(D_72), .O(ED_326) );
and2 gate( .a(CONST0), .b(D_72), .O(ED_327) );
and2 gate( .a(ED_324), .b(D_73_NOT), .O(ED_333) );
and2 gate( .a(ED_325), .b(D_73), .O(ED_331) );
and2 gate( .a(ED_326), .b(D_73_NOT), .O(ED_329) );
and2 gate( .a(ED_327), .b(D_73), .O(ED_328) );
or2  gate( .a(ED_328), .b(ED_329), .O(ED_330) );
or2  gate( .a(ED_330), .b(ED_331), .O(ED_332) );
or2  gate( .a(ED_333), .b(ED_332), .O(N422_OBF);
inv1 gate( .a(D_74), .O(D_74_NOT) );
inv1 gate( .a(D_75), .O(D_75_NOT) );
inv1 gate( .a(N425), .O(N425_NOT) );
and2 gate( .a(N425), .b(D_74_NOT), .O(ED_333) );
and2 gate( .a(N425_NOT), .b(D_74_NOT), .O(ED_334) );
and2 gate( .a(CONST1), .b(D_74), .O(ED_335) );
and2 gate( .a(CONST0), .b(D_74), .O(ED_336) );
and2 gate( .a(ED_333), .b(D_75_NOT), .O(ED_342) );
and2 gate( .a(ED_334), .b(D_75), .O(ED_340) );
and2 gate( .a(ED_335), .b(D_75_NOT), .O(ED_338) );
and2 gate( .a(ED_336), .b(D_75), .O(ED_337) );
or2  gate( .a(ED_337), .b(ED_338), .O(ED_339) );
or2  gate( .a(ED_339), .b(ED_340), .O(ED_341) );
or2  gate( .a(ED_342), .b(ED_341), .O(N425_OBF);
inv1 gate( .a(D_76), .O(D_76_NOT) );
inv1 gate( .a(D_77), .O(D_77_NOT) );
inv1 gate( .a(N429), .O(N429_NOT) );
and2 gate( .a(N429), .b(D_76_NOT), .O(ED_342) );
and2 gate( .a(N429_NOT), .b(D_76_NOT), .O(ED_343) );
and2 gate( .a(CONST1), .b(D_76), .O(ED_344) );
and2 gate( .a(CONST0), .b(D_76), .O(ED_345) );
and2 gate( .a(ED_342), .b(D_77_NOT), .O(ED_351) );
and2 gate( .a(ED_343), .b(D_77), .O(ED_349) );
and2 gate( .a(ED_344), .b(D_77_NOT), .O(ED_347) );
and2 gate( .a(ED_345), .b(D_77), .O(ED_346) );
or2  gate( .a(ED_346), .b(ED_347), .O(ED_348) );
or2  gate( .a(ED_348), .b(ED_349), .O(ED_350) );
or2  gate( .a(ED_351), .b(ED_350), .O(N429_OBF);
inv1 gate( .a(D_78), .O(D_78_NOT) );
inv1 gate( .a(D_79), .O(D_79_NOT) );
inv1 gate( .a(N432), .O(N432_NOT) );
and2 gate( .a(N432), .b(D_78_NOT), .O(ED_351) );
and2 gate( .a(N432_NOT), .b(D_78_NOT), .O(ED_352) );
and2 gate( .a(CONST1), .b(D_78), .O(ED_353) );
and2 gate( .a(CONST0), .b(D_78), .O(ED_354) );
and2 gate( .a(ED_351), .b(D_79_NOT), .O(ED_360) );
and2 gate( .a(ED_352), .b(D_79), .O(ED_358) );
and2 gate( .a(ED_353), .b(D_79_NOT), .O(ED_356) );
and2 gate( .a(ED_354), .b(D_79), .O(ED_355) );
or2  gate( .a(ED_355), .b(ED_356), .O(ED_357) );
or2  gate( .a(ED_357), .b(ED_358), .O(ED_359) );
or2  gate( .a(ED_360), .b(ED_359), .O(N432_OBF);
inv1 gate( .a(D_80), .O(D_80_NOT) );
inv1 gate( .a(D_81), .O(D_81_NOT) );
inv1 gate( .a(N381), .O(N381_NOT) );
and2 gate( .a(N381), .b(D_80_NOT), .O(ED_360) );
and2 gate( .a(N381_NOT), .b(D_80_NOT), .O(ED_361) );
and2 gate( .a(CONST1), .b(D_80), .O(ED_362) );
and2 gate( .a(CONST0), .b(D_80), .O(ED_363) );
and2 gate( .a(ED_360), .b(D_81_NOT), .O(ED_369) );
and2 gate( .a(ED_361), .b(D_81), .O(ED_367) );
and2 gate( .a(ED_362), .b(D_81_NOT), .O(ED_365) );
and2 gate( .a(ED_363), .b(D_81), .O(ED_364) );
or2  gate( .a(ED_364), .b(ED_365), .O(ED_366) );
or2  gate( .a(ED_366), .b(ED_367), .O(ED_368) );
or2  gate( .a(ED_369), .b(ED_368), .O(N381_OBF);
inv1 gate( .a(D_82), .O(D_82_NOT) );
inv1 gate( .a(D_83), .O(D_83_NOT) );
inv1 gate( .a(N386), .O(N386_NOT) );
and2 gate( .a(N386), .b(D_82_NOT), .O(ED_369) );
and2 gate( .a(N386_NOT), .b(D_82_NOT), .O(ED_370) );
and2 gate( .a(CONST1), .b(D_82), .O(ED_371) );
and2 gate( .a(CONST0), .b(D_82), .O(ED_372) );
and2 gate( .a(ED_369), .b(D_83_NOT), .O(ED_378) );
and2 gate( .a(ED_370), .b(D_83), .O(ED_376) );
and2 gate( .a(ED_371), .b(D_83_NOT), .O(ED_374) );
and2 gate( .a(ED_372), .b(D_83), .O(ED_373) );
or2  gate( .a(ED_373), .b(ED_374), .O(ED_375) );
or2  gate( .a(ED_375), .b(ED_376), .O(ED_377) );
or2  gate( .a(ED_378), .b(ED_377), .O(N386_OBF);
inv1 gate( .a(D_84), .O(D_84_NOT) );
inv1 gate( .a(D_85), .O(D_85_NOT) );
inv1 gate( .a(N425), .O(N425_NOT) );
and2 gate( .a(N425), .b(D_84_NOT), .O(ED_378) );
and2 gate( .a(N425_NOT), .b(D_84_NOT), .O(ED_379) );
and2 gate( .a(CONST1), .b(D_84), .O(ED_380) );
and2 gate( .a(CONST0), .b(D_84), .O(ED_381) );
and2 gate( .a(ED_378), .b(D_85_NOT), .O(ED_387) );
and2 gate( .a(ED_379), .b(D_85), .O(ED_385) );
and2 gate( .a(ED_380), .b(D_85_NOT), .O(ED_383) );
and2 gate( .a(ED_381), .b(D_85), .O(ED_382) );
or2  gate( .a(ED_382), .b(ED_383), .O(ED_384) );
or2  gate( .a(ED_384), .b(ED_385), .O(ED_386) );
or2  gate( .a(ED_387), .b(ED_386), .O(N425_OBF);
inv1 gate( .a(D_86), .O(D_86_NOT) );
inv1 gate( .a(D_87), .O(D_87_NOT) );
inv1 gate( .a(N428), .O(N428_NOT) );
and2 gate( .a(N428), .b(D_86_NOT), .O(ED_387) );
and2 gate( .a(N428_NOT), .b(D_86_NOT), .O(ED_388) );
and2 gate( .a(CONST1), .b(D_86), .O(ED_389) );
and2 gate( .a(CONST0), .b(D_86), .O(ED_390) );
and2 gate( .a(ED_387), .b(D_87_NOT), .O(ED_396) );
and2 gate( .a(ED_388), .b(D_87), .O(ED_394) );
and2 gate( .a(ED_389), .b(D_87_NOT), .O(ED_392) );
and2 gate( .a(ED_390), .b(D_87), .O(ED_391) );
or2  gate( .a(ED_391), .b(ED_392), .O(ED_393) );
or2  gate( .a(ED_393), .b(ED_394), .O(ED_395) );
or2  gate( .a(ED_396), .b(ED_395), .O(N428_OBF);
inv1 gate( .a(D_88), .O(D_88_NOT) );
inv1 gate( .a(D_89), .O(D_89_NOT) );
inv1 gate( .a(N431), .O(N431_NOT) );
and2 gate( .a(N431), .b(D_88_NOT), .O(ED_396) );
and2 gate( .a(N431_NOT), .b(D_88_NOT), .O(ED_397) );
and2 gate( .a(CONST1), .b(D_88), .O(ED_398) );
and2 gate( .a(CONST0), .b(D_88), .O(ED_399) );
and2 gate( .a(ED_396), .b(D_89_NOT), .O(ED_405) );
and2 gate( .a(ED_397), .b(D_89), .O(ED_403) );
and2 gate( .a(ED_398), .b(D_89_NOT), .O(ED_401) );
and2 gate( .a(ED_399), .b(D_89), .O(ED_400) );
or2  gate( .a(ED_400), .b(ED_401), .O(ED_402) );
or2  gate( .a(ED_402), .b(ED_403), .O(ED_404) );
or2  gate( .a(ED_405), .b(ED_404), .O(N431_OBF);
inv1 gate( .a(D_90), .O(D_90_NOT) );
inv1 gate( .a(D_91), .O(D_91_NOT) );
inv1 gate( .a(N258), .O(N258_NOT) );
and2 gate( .a(N258), .b(D_90_NOT), .O(ED_405) );
and2 gate( .a(N258_NOT), .b(D_90_NOT), .O(ED_406) );
and2 gate( .a(CONST1), .b(D_90), .O(ED_407) );
and2 gate( .a(CONST0), .b(D_90), .O(ED_408) );
and2 gate( .a(ED_405), .b(D_91_NOT), .O(ED_414) );
and2 gate( .a(ED_406), .b(D_91), .O(ED_412) );
and2 gate( .a(ED_407), .b(D_91_NOT), .O(ED_410) );
and2 gate( .a(ED_408), .b(D_91), .O(ED_409) );
or2  gate( .a(ED_409), .b(ED_410), .O(ED_411) );
or2  gate( .a(ED_411), .b(ED_412), .O(ED_413) );
or2  gate( .a(ED_414), .b(ED_413), .O(N258_OBF);
inv1 gate( .a(D_92), .O(D_92_NOT) );
inv1 gate( .a(D_93), .O(D_93_NOT) );
inv1 gate( .a(N346), .O(N346_NOT) );
and2 gate( .a(N346), .b(D_92_NOT), .O(ED_414) );
and2 gate( .a(N346_NOT), .b(D_92_NOT), .O(ED_415) );
and2 gate( .a(CONST1), .b(D_92), .O(ED_416) );
and2 gate( .a(CONST0), .b(D_92), .O(ED_417) );
and2 gate( .a(ED_414), .b(D_93_NOT), .O(ED_423) );
and2 gate( .a(ED_415), .b(D_93), .O(ED_421) );
and2 gate( .a(ED_416), .b(D_93_NOT), .O(ED_419) );
and2 gate( .a(ED_417), .b(D_93), .O(ED_418) );
or2  gate( .a(ED_418), .b(ED_419), .O(ED_420) );
or2  gate( .a(ED_420), .b(ED_421), .O(ED_422) );
or2  gate( .a(ED_423), .b(ED_422), .O(N346_OBF);
inv1 gate( .a(D_94), .O(D_94_NOT) );
inv1 gate( .a(D_95), .O(D_95_NOT) );
inv1 gate( .a(N378), .O(N378_NOT) );
and2 gate( .a(N378), .b(D_94_NOT), .O(ED_423) );
and2 gate( .a(N378_NOT), .b(D_94_NOT), .O(ED_424) );
and2 gate( .a(CONST1), .b(D_94), .O(ED_425) );
and2 gate( .a(CONST0), .b(D_94), .O(ED_426) );
and2 gate( .a(ED_423), .b(D_95_NOT), .O(ED_432) );
and2 gate( .a(ED_424), .b(D_95), .O(ED_430) );
and2 gate( .a(ED_425), .b(D_95_NOT), .O(ED_428) );
and2 gate( .a(ED_426), .b(D_95), .O(ED_427) );
or2  gate( .a(ED_427), .b(ED_428), .O(ED_429) );
or2  gate( .a(ED_429), .b(ED_430), .O(ED_431) );
or2  gate( .a(ED_432), .b(ED_431), .O(N378_OBF);
inv1 gate( .a(D_96), .O(D_96_NOT) );
inv1 gate( .a(D_97), .O(D_97_NOT) );
inv1 gate( .a(N95), .O(N95_NOT) );
and2 gate( .a(N95), .b(D_96_NOT), .O(ED_432) );
and2 gate( .a(N95_NOT), .b(D_96_NOT), .O(ED_433) );
and2 gate( .a(CONST1), .b(D_96), .O(ED_434) );
and2 gate( .a(CONST0), .b(D_96), .O(ED_435) );
and2 gate( .a(ED_432), .b(D_97_NOT), .O(ED_441) );
and2 gate( .a(ED_433), .b(D_97), .O(ED_439) );
and2 gate( .a(ED_434), .b(D_97_NOT), .O(ED_437) );
and2 gate( .a(ED_435), .b(D_97), .O(ED_436) );
or2  gate( .a(ED_436), .b(ED_437), .O(ED_438) );
or2  gate( .a(ED_438), .b(ED_439), .O(ED_440) );
or2  gate( .a(ED_441), .b(ED_440), .O(N95_OBF);
inv1 gate( .a(D_98), .O(D_98_NOT) );
inv1 gate( .a(D_99), .O(D_99_NOT) );
inv1 gate( .a(N411), .O(N411_NOT) );
and2 gate( .a(N411), .b(D_98_NOT), .O(ED_441) );
and2 gate( .a(N411_NOT), .b(D_98_NOT), .O(ED_442) );
and2 gate( .a(CONST1), .b(D_98), .O(ED_443) );
and2 gate( .a(CONST0), .b(D_98), .O(ED_444) );
and2 gate( .a(ED_441), .b(D_99_NOT), .O(ED_450) );
and2 gate( .a(ED_442), .b(D_99), .O(ED_448) );
and2 gate( .a(ED_443), .b(D_99_NOT), .O(ED_446) );
and2 gate( .a(ED_444), .b(D_99), .O(ED_445) );
or2  gate( .a(ED_445), .b(ED_446), .O(ED_447) );
or2  gate( .a(ED_447), .b(ED_448), .O(ED_449) );
or2  gate( .a(ED_450), .b(ED_449), .O(N411_OBF);

endmodule
